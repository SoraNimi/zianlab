** Generated for: hspiceD
** Generated on: Jun 13 21:33:30 2018
** Design library name: reram
** Design cell name: XORNET4
** Design view name: schematic
.PARAM blinresistor=2000
.PARAM blresistor=3000

.TRAN 10e-12 200e-9 START=0.0

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.OPTION PROBE=1

.PROBE tran v(l0bl0)
.PROBE tran v(l0bl1)
.PROBE tran v(l0bl2)
.PROBE tran v(l0bl3)
.PROBE tran v(l0bl4)
.PROBE tran v(l0bl5)
.PROBE tran v(l0bl6)
.PROBE tran v(l0bl7)
.PROBE tran v(l0bl8)
.PROBE tran v(l0bl9)
.PROBE tran v(l0bl10)
.PROBE tran v(l0bl11)
.PROBE tran v(l0bl12)
.PROBE tran v(l0bl13)
.PROBE tran v(l0bl14)
.PROBE tran v(l0bl15)
.PROBE tran v(l0bl16)
.PROBE tran v(l0bl17)
.PROBE tran v(l0bl18)
.PROBE tran v(l0bl19)
.PROBE tran v(l0bl20)
.PROBE tran v(l0bl21)
.PROBE tran v(l0bl22)
.PROBE tran v(l0bl23)
.PROBE tran v(l0bl24)
.PROBE tran v(l0bl25)
.PROBE tran v(l0bl26)
.PROBE tran v(l0bl27)
.PROBE tran v(l0bl28)
.PROBE tran v(l0bl29)
.PROBE tran v(l0bl30)
.PROBE tran v(l0bl31)
.PROBE tran v(l0bl32)
.PROBE tran v(l0bl33)
.PROBE tran v(l0bl34)
.PROBE tran v(l0bl35)
.PROBE tran v(l0bl36)
.PROBE tran v(l0bl37)
.PROBE tran v(l0bl38)
.PROBE tran v(l0bl39)
.PROBE tran v(l0bl40)
.PROBE tran v(l0bl41)
.PROBE tran v(l0bl42)
.PROBE tran v(l0bl43)
.PROBE tran v(l0bl44)
.PROBE tran v(l0bl45)
.PROBE tran v(l0bl46)
.PROBE tran v(l0bl47)
.PROBE tran v(l0bl48)
.PROBE tran v(l0bl49)
.PROBE tran v(l0bl50)
.PROBE tran v(l0bl51)
.PROBE tran v(l0bl52)
.PROBE tran v(l0bl53)
.PROBE tran v(l0bl54)
.PROBE tran v(l0bl55)
.PROBE tran v(l0bl56)
.PROBE tran v(l0bl57)
.PROBE tran v(l0bl58)
.PROBE tran v(l0bl59)
.PROBE tran v(l0bl60)
.PROBE tran v(l0bl61)
.PROBE tran v(l0bl62)
.PROBE tran v(l0bl63)
.PROBE tran v(l0bl64)
.PROBE tran v(l0bl65)
.PROBE tran v(l0bl66)
.PROBE tran v(l0bl67)
.PROBE tran v(l0bl68)
.PROBE tran v(l0bl69)
.PROBE tran v(l0bl70)
.PROBE tran v(l0bl71)
.PROBE tran v(l0bl72)
.PROBE tran v(l0bl73)
.PROBE tran v(l0bl74)
.PROBE tran v(l0bl75)
.PROBE tran v(l0bl76)
.PROBE tran v(l0bl77)
.PROBE tran v(l0bl78)
.PROBE tran v(l0bl79)
.PROBE tran v(l0bl80)
.PROBE tran v(l0bl81)
.PROBE tran v(l0bl82)
.PROBE tran v(l0bl83)
.PROBE tran v(l0bl84)
.PROBE tran v(l0bl85)
.PROBE tran v(l0bl86)
.PROBE tran v(l0bl87)
.PROBE tran v(l0bl88)
.PROBE tran v(l0bl89)
.PROBE tran v(l0bl90)
.PROBE tran v(l0bl91)
.PROBE tran v(l0bl92)
.PROBE tran v(l0bl93)
.PROBE tran v(l0bl94)
.PROBE tran v(l0bl95)
.PROBE tran v(l0bl96)
.PROBE tran v(l0bl97)
.PROBE tran v(l0bl98)
.PROBE tran v(l0bl99)
.PROBE tran v(l0bl100)
.PROBE tran v(l0bl101)
.PROBE tran v(l0bl102)
.PROBE tran v(l0bl103)
.PROBE tran v(l0bl104)
.PROBE tran v(l0bl105)
.PROBE tran v(l0bl106)
.PROBE tran v(l0bl107)
.PROBE tran v(l0bl108)
.PROBE tran v(l0bl109)
.PROBE tran v(l0bl110)
.PROBE tran v(l0bl111)
.PROBE tran v(l0bl112)
.PROBE tran v(l0bl113)
.PROBE tran v(l0bl114)
.PROBE tran v(l0bl115)
.PROBE tran v(l0bl116)
.PROBE tran v(l0bl117)
.PROBE tran v(l0bl118)
.PROBE tran v(l0bl119)
.PROBE tran v(l0bl120)
.PROBE tran v(l0bl121)
.PROBE tran v(l0bl122)
.PROBE tran v(l0bl123)
.PROBE tran v(l0bl124)
.PROBE tran v(l0bl125)
.PROBE tran v(l0bl126)
.PROBE tran v(l0bl127)
.PROBE tran v(l0bl128)
.PROBE tran v(l0bl129)
.PROBE tran v(l0bl130)
.PROBE tran v(l0bl131)
.PROBE tran v(l0bl132)
.PROBE tran v(l0bl133)
.PROBE tran v(l0bl134)
.PROBE tran v(l0bl135)
.PROBE tran v(l0bl136)
.PROBE tran v(l0bl137)
.PROBE tran v(l0bl138)
.PROBE tran v(l0bl139)
.PROBE tran v(l0bl140)
.PROBE tran v(l0bl141)
.PROBE tran v(l0bl142)
.PROBE tran v(l0bl143)
.PROBE tran v(l0bl144)
.PROBE tran v(l0bl145)
.PROBE tran v(l0bl146)
.PROBE tran v(l0bl147)
.PROBE tran v(l0bl148)
.PROBE tran v(l0bl149)
.PROBE tran v(l0bl150)
.PROBE tran v(l0bl151)
.PROBE tran v(l0bl152)
.PROBE tran v(l0bl153)
.PROBE tran v(l0bl154)
.PROBE tran v(l0bl155)
.PROBE tran v(l0bl156)
.PROBE tran v(l0bl157)
.PROBE tran v(l0bl158)
.PROBE tran v(l0bl159)
.PROBE tran v(l0bl160)
.PROBE tran v(l0bl161)
.PROBE tran v(l0bl162)
.PROBE tran v(l0bl163)
.PROBE tran v(l0bl164)
.PROBE tran v(l0bl165)
.PROBE tran v(l0bl166)
.PROBE tran v(l0bl167)
.PROBE tran v(l0bl168)
.PROBE tran v(l0bl169)
.PROBE tran v(l0bl170)
.PROBE tran v(l0bl171)
.PROBE tran v(l0bl172)
.PROBE tran v(l0bl173)
.PROBE tran v(l0bl174)
.PROBE tran v(l0bl175)
.PROBE tran v(l0bl176)
.PROBE tran v(l0bl177)
.PROBE tran v(l0bl178)
.PROBE tran v(l0bl179)
.PROBE tran v(l0bl180)
.PROBE tran v(l0bl181)
.PROBE tran v(l0bl182)
.PROBE tran v(l0bl183)
.PROBE tran v(l0bl184)
.PROBE tran v(l0bl185)
.PROBE tran v(l0bl186)
.PROBE tran v(l0bl187)
.PROBE tran v(l0bl188)
.PROBE tran v(l0bl189)
.PROBE tran v(l0bl190)
.PROBE tran v(l0bl191)
.PROBE tran v(l0bl192)
.PROBE tran v(l0bl193)
.PROBE tran v(l0bl194)
.PROBE tran v(l0bl195)
.PROBE tran v(l0bl196)
.PROBE tran v(l0bl197)
.PROBE tran v(l0bl198)
.PROBE tran v(l0bl199)
.PROBE tran v(l0bl200)
.PROBE tran v(l0bl201)
.PROBE tran v(l0bl202)
.PROBE tran v(l0bl203)
.PROBE tran v(l0bl204)
.PROBE tran v(l0bl205)
.PROBE tran v(l0bl206)
.PROBE tran v(l0bl207)
.PROBE tran v(l0bl208)
.PROBE tran v(l0bl209)
.PROBE tran v(l0bl210)
.PROBE tran v(l0bl211)
.PROBE tran v(l0bl212)
.PROBE tran v(l0bl213)
.PROBE tran v(l0bl214)
.PROBE tran v(l0bl215)
.PROBE tran v(l0bl216)
.PROBE tran v(l0bl217)
.PROBE tran v(l0bl218)
.PROBE tran v(l0bl219)
.PROBE tran v(l0bl220)
.PROBE tran v(l0bl221)
.PROBE tran v(l0bl222)
.PROBE tran v(l0bl223)
.PROBE tran v(l0bl224)
.PROBE tran v(l0bl225)
.PROBE tran v(l0bl226)
.PROBE tran v(l0bl227)
.PROBE tran v(l0bl228)
.PROBE tran v(l0bl229)
.PROBE tran v(l0bl230)
.PROBE tran v(l0bl231)
.PROBE tran v(l0bl232)
.PROBE tran v(l0bl233)
.PROBE tran v(l0bl234)
.PROBE tran v(l0bl235)
.PROBE tran v(l0bl236)
.PROBE tran v(l0bl237)
.PROBE tran v(l0bl238)
.PROBE tran v(l0bl239)
.PROBE tran v(l0bl240)
.PROBE tran v(l0bl241)
.PROBE tran v(l0bl242)
.PROBE tran v(l0bl243)
.PROBE tran v(l0bl244)
.PROBE tran v(l0bl245)
.PROBE tran v(l0bl246)
.PROBE tran v(l0bl247)
.PROBE tran v(l0bl248)
.PROBE tran v(l0bl249)
.PROBE tran v(l0bl250)
.PROBE tran v(l0bl251)
.PROBE tran v(l0bl252)
.PROBE tran v(l0bl253)
.PROBE tran v(l0bl254)
.PROBE tran v(l0bl255)
.PROBE tran v(l0bl256)
.PROBE tran v(l0bl257)
.PROBE tran v(l0bl258)
.PROBE tran v(l0bl259)
.PROBE tran v(l0bl260)
.PROBE tran v(l0bl261)
.PROBE tran v(l0bl262)
.PROBE tran v(l0bl263)
.PROBE tran v(l0bl264)
.PROBE tran v(l0bl265)
.PROBE tran v(l0bl266)
.PROBE tran v(l0bl267)
.PROBE tran v(l0bl268)
.PROBE tran v(l0bl269)
.PROBE tran v(l0bl270)
.PROBE tran v(l0bl271)
.PROBE tran v(l0bl272)
.PROBE tran v(l0bl273)
.PROBE tran v(l0bl274)
.PROBE tran v(l0bl275)
.PROBE tran v(l0bl276)
.PROBE tran v(l0bl277)
.PROBE tran v(l0bl278)
.PROBE tran v(l0bl279)
.PROBE tran v(l0bl280)
.PROBE tran v(l0bl281)
.PROBE tran v(l0bl282)
.PROBE tran v(l0bl283)
.PROBE tran v(l0bl284)
.PROBE tran v(l0bl285)
.PROBE tran v(l0bl286)
.PROBE tran v(l0bl287)
.PROBE tran v(l0bl288)
.PROBE tran v(l0bl289)
.PROBE tran v(l0bl290)
.PROBE tran v(l0bl291)
.PROBE tran v(l0bl292)
.PROBE tran v(l0bl293)
.PROBE tran v(l0bl294)
.PROBE tran v(l0bl295)
.PROBE tran v(l0bl296)
.PROBE tran v(l0bl297)
.PROBE tran v(l0bl298)
.PROBE tran v(l0bl299)
.PROBE tran v(l0bl300)
.PROBE tran v(l0bl301)
.PROBE tran v(l0bl302)
.PROBE tran v(l0bl303)
.PROBE tran v(l0bl304)
.PROBE tran v(l0bl305)
.PROBE tran v(l0bl306)
.PROBE tran v(l0bl307)
.PROBE tran v(l0bl308)
.PROBE tran v(l0bl309)
.PROBE tran v(l0bl310)
.PROBE tran v(l0bl311)
.PROBE tran v(l0bl312)
.PROBE tran v(l0bl313)
.PROBE tran v(l0bl314)
.PROBE tran v(l0bl315)
.PROBE tran v(l0bl316)
.PROBE tran v(l0bl317)
.PROBE tran v(l0bl318)
.PROBE tran v(l0bl319)
.PROBE tran v(l0bl320)
.PROBE tran v(l0bl321)
.PROBE tran v(l0bl322)
.PROBE tran v(l0bl323)
.PROBE tran v(l0bl324)
.PROBE tran v(l0bl325)
.PROBE tran v(l0bl326)
.PROBE tran v(l0bl327)
.PROBE tran v(l0bl328)
.PROBE tran v(l0bl329)
.PROBE tran v(l0bl330)
.PROBE tran v(l0bl331)
.PROBE tran v(l0bl332)
.PROBE tran v(l0bl333)
.PROBE tran v(l0bl334)
.PROBE tran v(l0bl335)
.PROBE tran v(l0bl336)
.PROBE tran v(l0bl337)
.PROBE tran v(l0bl338)
.PROBE tran v(l0bl339)
.PROBE tran v(l0bl340)
.PROBE tran v(l0bl341)
.PROBE tran v(l0bl342)
.PROBE tran v(l0bl343)
.PROBE tran v(l0bl344)
.PROBE tran v(l0bl345)
.PROBE tran v(l0bl346)
.PROBE tran v(l0bl347)
.PROBE tran v(l0bl348)
.PROBE tran v(l0bl349)
.PROBE tran v(l0bl350)
.PROBE tran v(l0bl351)
.PROBE tran v(l0bl352)
.PROBE tran v(l0bl353)
.PROBE tran v(l0bl354)
.PROBE tran v(l0bl355)
.PROBE tran v(l0bl356)
.PROBE tran v(l0bl357)
.PROBE tran v(l0bl358)
.PROBE tran v(l0bl359)
.PROBE tran v(l0bl360)
.PROBE tran v(l0bl361)
.PROBE tran v(l0bl362)
.PROBE tran v(l0bl363)
.PROBE tran v(l0bl364)
.PROBE tran v(l0bl365)
.PROBE tran v(l0bl366)
.PROBE tran v(l0bl367)
.PROBE tran v(l0bl368)
.PROBE tran v(l0bl369)
.PROBE tran v(l0bl370)
.PROBE tran v(l0bl371)
.PROBE tran v(l0bl372)
.PROBE tran v(l0bl373)
.PROBE tran v(l0bl374)
.PROBE tran v(l0bl375)
.PROBE tran v(l0bl376)
.PROBE tran v(l0bl377)
.PROBE tran v(l0bl378)
.PROBE tran v(l0bl379)
.PROBE tran v(l0bl380)
.PROBE tran v(l0bl381)
.PROBE tran v(l0bl382)
.PROBE tran v(l0bl383)
.PROBE tran v(l0bl384)
.PROBE tran v(l0bl385)
.PROBE tran v(l0bl386)
.PROBE tran v(l0bl387)
.PROBE tran v(l0bl388)
.PROBE tran v(l0bl389)
.PROBE tran v(l0bl390)
.PROBE tran v(l0bl391)
.PROBE tran v(l0bl392)
.PROBE tran v(l0bl393)
.PROBE tran v(l0bl394)
.PROBE tran v(l0bl395)
.PROBE tran v(l0bl396)
.PROBE tran v(l0bl397)
.PROBE tran v(l0bl398)
.PROBE tran v(l0bl399)
.PROBE tran v(l0bl400)
.PROBE tran v(l0bl401)
.PROBE tran v(l0bl402)
.PROBE tran v(l0bl403)
.PROBE tran v(l0bl404)
.PROBE tran v(l0bl405)
.PROBE tran v(l0bl406)
.PROBE tran v(l0bl407)
.PROBE tran v(l0bl408)
.PROBE tran v(l0bl409)
.PROBE tran v(l0bl410)
.PROBE tran v(l0bl411)
.PROBE tran v(l0bl412)
.PROBE tran v(l0bl413)
.PROBE tran v(l0bl414)
.PROBE tran v(l0bl415)
.PROBE tran v(l0bl416)
.PROBE tran v(l0bl417)
.PROBE tran v(l0bl418)
.PROBE tran v(l0bl419)
.PROBE tran v(l0bl420)
.PROBE tran v(l0bl421)
.PROBE tran v(l0bl422)
.PROBE tran v(l0bl423)
.PROBE tran v(l0bl424)
.PROBE tran v(l0bl425)
.PROBE tran v(l0bl426)
.PROBE tran v(l0bl427)
.PROBE tran v(l0bl428)
.PROBE tran v(l0bl429)
.PROBE tran v(l0bl430)
.PROBE tran v(l0bl431)
.PROBE tran v(l0bl432)
.PROBE tran v(l0bl433)
.PROBE tran v(l0bl434)
.PROBE tran v(l0bl435)
.PROBE tran v(l0bl436)
.PROBE tran v(l0bl437)
.PROBE tran v(l0bl438)
.PROBE tran v(l0bl439)
.PROBE tran v(l0bl440)
.PROBE tran v(l0bl441)
.PROBE tran v(l0bl442)
.PROBE tran v(l0bl443)
.PROBE tran v(l0bl444)
.PROBE tran v(l0bl445)
.PROBE tran v(l0bl446)
.PROBE tran v(l0bl447)
.PROBE tran v(l0bl448)
.PROBE tran v(l0bl449)
.PROBE tran v(l0bl450)
.PROBE tran v(l0bl451)
.PROBE tran v(l0bl452)
.PROBE tran v(l0bl453)
.PROBE tran v(l0bl454)
.PROBE tran v(l0bl455)
.PROBE tran v(l0bl456)
.PROBE tran v(l0bl457)
.PROBE tran v(l0bl458)
.PROBE tran v(l0bl459)
.PROBE tran v(l0bl460)
.PROBE tran v(l0bl461)
.PROBE tran v(l0bl462)
.PROBE tran v(l0bl463)
.PROBE tran v(l0bl464)
.PROBE tran v(l0bl465)
.PROBE tran v(l0bl466)
.PROBE tran v(l0bl467)
.PROBE tran v(l0bl468)
.PROBE tran v(l0bl469)
.PROBE tran v(l0bl470)
.PROBE tran v(l0bl471)
.PROBE tran v(l0bl472)
.PROBE tran v(l0bl473)
.PROBE tran v(l0bl474)
.PROBE tran v(l0bl475)
.PROBE tran v(l0bl476)
.PROBE tran v(l0bl477)
.PROBE tran v(l0bl478)
.PROBE tran v(l0bl479)
.PROBE tran v(l0bl480)
.PROBE tran v(l0bl481)
.PROBE tran v(l0bl482)
.PROBE tran v(l0bl483)
.PROBE tran v(l0bl484)
.PROBE tran v(l0bl485)
.PROBE tran v(l0bl486)
.PROBE tran v(l0bl487)
.PROBE tran v(l0bl488)
.PROBE tran v(l0bl489)
.PROBE tran v(l0bl490)
.PROBE tran v(l0bl491)
.PROBE tran v(l0bl492)
.PROBE tran v(l0bl493)
.PROBE tran v(l0bl494)
.PROBE tran v(l0bl495)
.PROBE tran v(l0bl496)
.PROBE tran v(l0bl497)
.PROBE tran v(l0bl498)
.PROBE tran v(l0bl499)
.PROBE tran v(l0bl500)
.PROBE tran v(l0bl501)
.PROBE tran v(l0bl502)
.PROBE tran v(l0bl503)
.PROBE tran v(l0bl504)
.PROBE tran v(l0bl505)
.PROBE tran v(l0bl506)
.PROBE tran v(l0bl507)
.PROBE tran v(l0bl508)
.PROBE tran v(l0bl509)
.PROBE tran v(l0bl510)
.PROBE tran v(l0bl511)

.PROBE tran v(l1bl0)
.PROBE tran v(l1bl1)
.PROBE tran v(l1bl2)
.PROBE tran v(l1bl3)
.PROBE tran v(l1bl4)
.PROBE tran v(l1bl5)
.PROBE tran v(l1bl6)
.PROBE tran v(l1bl7)
.PROBE tran v(l1bl8)
.PROBE tran v(l1bl9)
.PROBE tran v(l1bl10)
.PROBE tran v(l1bl11)
.PROBE tran v(l1bl12)
.PROBE tran v(l1bl13)
.PROBE tran v(l1bl14)
.PROBE tran v(l1bl15)
.PROBE tran v(l1bl16)
.PROBE tran v(l1bl17)
.PROBE tran v(l1bl18)
.PROBE tran v(l1bl19)
.PROBE tran v(l1bl20)
.PROBE tran v(l1bl21)
.PROBE tran v(l1bl22)
.PROBE tran v(l1bl23)
.PROBE tran v(l1bl24)
.PROBE tran v(l1bl25)
.PROBE tran v(l1bl26)
.PROBE tran v(l1bl27)
.PROBE tran v(l1bl28)
.PROBE tran v(l1bl29)
.PROBE tran v(l1bl30)
.PROBE tran v(l1bl31)
.PROBE tran v(l1bl32)
.PROBE tran v(l1bl33)
.PROBE tran v(l1bl34)
.PROBE tran v(l1bl35)
.PROBE tran v(l1bl36)
.PROBE tran v(l1bl37)
.PROBE tran v(l1bl38)
.PROBE tran v(l1bl39)
.PROBE tran v(l1bl40)
.PROBE tran v(l1bl41)
.PROBE tran v(l1bl42)
.PROBE tran v(l1bl43)
.PROBE tran v(l1bl44)
.PROBE tran v(l1bl45)
.PROBE tran v(l1bl46)
.PROBE tran v(l1bl47)
.PROBE tran v(l1bl48)
.PROBE tran v(l1bl49)
.PROBE tran v(l1bl50)
.PROBE tran v(l1bl51)
.PROBE tran v(l1bl52)
.PROBE tran v(l1bl53)
.PROBE tran v(l1bl54)
.PROBE tran v(l1bl55)
.PROBE tran v(l1bl56)
.PROBE tran v(l1bl57)
.PROBE tran v(l1bl58)
.PROBE tran v(l1bl59)
.PROBE tran v(l1bl60)
.PROBE tran v(l1bl61)
.PROBE tran v(l1bl62)
.PROBE tran v(l1bl63)
.PROBE tran v(l1bl64)
.PROBE tran v(l1bl65)
.PROBE tran v(l1bl66)
.PROBE tran v(l1bl67)
.PROBE tran v(l1bl68)
.PROBE tran v(l1bl69)
.PROBE tran v(l1bl70)
.PROBE tran v(l1bl71)
.PROBE tran v(l1bl72)
.PROBE tran v(l1bl73)
.PROBE tran v(l1bl74)
.PROBE tran v(l1bl75)
.PROBE tran v(l1bl76)
.PROBE tran v(l1bl77)
.PROBE tran v(l1bl78)
.PROBE tran v(l1bl79)
.PROBE tran v(l1bl80)
.PROBE tran v(l1bl81)
.PROBE tran v(l1bl82)
.PROBE tran v(l1bl83)
.PROBE tran v(l1bl84)
.PROBE tran v(l1bl85)
.PROBE tran v(l1bl86)
.PROBE tran v(l1bl87)
.PROBE tran v(l1bl88)
.PROBE tran v(l1bl89)
.PROBE tran v(l1bl90)
.PROBE tran v(l1bl91)
.PROBE tran v(l1bl92)
.PROBE tran v(l1bl93)
.PROBE tran v(l1bl94)
.PROBE tran v(l1bl95)
.PROBE tran v(l1bl96)
.PROBE tran v(l1bl97)
.PROBE tran v(l1bl98)
.PROBE tran v(l1bl99)
.PROBE tran v(l1bl100)
.PROBE tran v(l1bl101)
.PROBE tran v(l1bl102)
.PROBE tran v(l1bl103)
.PROBE tran v(l1bl104)
.PROBE tran v(l1bl105)
.PROBE tran v(l1bl106)
.PROBE tran v(l1bl107)
.PROBE tran v(l1bl108)
.PROBE tran v(l1bl109)
.PROBE tran v(l1bl110)
.PROBE tran v(l1bl111)
.PROBE tran v(l1bl112)
.PROBE tran v(l1bl113)
.PROBE tran v(l1bl114)
.PROBE tran v(l1bl115)
.PROBE tran v(l1bl116)
.PROBE tran v(l1bl117)
.PROBE tran v(l1bl118)
.PROBE tran v(l1bl119)
.PROBE tran v(l1bl120)
.PROBE tran v(l1bl121)
.PROBE tran v(l1bl122)
.PROBE tran v(l1bl123)
.PROBE tran v(l1bl124)
.PROBE tran v(l1bl125)
.PROBE tran v(l1bl126)
.PROBE tran v(l1bl127)
.PROBE tran v(l1bl128)
.PROBE tran v(l1bl129)
.PROBE tran v(l1bl130)
.PROBE tran v(l1bl131)
.PROBE tran v(l1bl132)
.PROBE tran v(l1bl133)
.PROBE tran v(l1bl134)
.PROBE tran v(l1bl135)
.PROBE tran v(l1bl136)
.PROBE tran v(l1bl137)
.PROBE tran v(l1bl138)
.PROBE tran v(l1bl139)
.PROBE tran v(l1bl140)
.PROBE tran v(l1bl141)
.PROBE tran v(l1bl142)
.PROBE tran v(l1bl143)
.PROBE tran v(l1bl144)
.PROBE tran v(l1bl145)
.PROBE tran v(l1bl146)
.PROBE tran v(l1bl147)
.PROBE tran v(l1bl148)
.PROBE tran v(l1bl149)
.PROBE tran v(l1bl150)
.PROBE tran v(l1bl151)
.PROBE tran v(l1bl152)
.PROBE tran v(l1bl153)
.PROBE tran v(l1bl154)
.PROBE tran v(l1bl155)
.PROBE tran v(l1bl156)
.PROBE tran v(l1bl157)
.PROBE tran v(l1bl158)
.PROBE tran v(l1bl159)
.PROBE tran v(l1bl160)
.PROBE tran v(l1bl161)
.PROBE tran v(l1bl162)
.PROBE tran v(l1bl163)
.PROBE tran v(l1bl164)
.PROBE tran v(l1bl165)
.PROBE tran v(l1bl166)
.PROBE tran v(l1bl167)
.PROBE tran v(l1bl168)
.PROBE tran v(l1bl169)
.PROBE tran v(l1bl170)
.PROBE tran v(l1bl171)
.PROBE tran v(l1bl172)
.PROBE tran v(l1bl173)
.PROBE tran v(l1bl174)
.PROBE tran v(l1bl175)
.PROBE tran v(l1bl176)
.PROBE tran v(l1bl177)
.PROBE tran v(l1bl178)
.PROBE tran v(l1bl179)
.PROBE tran v(l1bl180)
.PROBE tran v(l1bl181)
.PROBE tran v(l1bl182)
.PROBE tran v(l1bl183)
.PROBE tran v(l1bl184)
.PROBE tran v(l1bl185)
.PROBE tran v(l1bl186)
.PROBE tran v(l1bl187)
.PROBE tran v(l1bl188)
.PROBE tran v(l1bl189)
.PROBE tran v(l1bl190)
.PROBE tran v(l1bl191)
.PROBE tran v(l1bl192)
.PROBE tran v(l1bl193)
.PROBE tran v(l1bl194)
.PROBE tran v(l1bl195)
.PROBE tran v(l1bl196)
.PROBE tran v(l1bl197)
.PROBE tran v(l1bl198)
.PROBE tran v(l1bl199)
.PROBE tran v(l1bl200)
.PROBE tran v(l1bl201)
.PROBE tran v(l1bl202)
.PROBE tran v(l1bl203)
.PROBE tran v(l1bl204)
.PROBE tran v(l1bl205)
.PROBE tran v(l1bl206)
.PROBE tran v(l1bl207)
.PROBE tran v(l1bl208)
.PROBE tran v(l1bl209)
.PROBE tran v(l1bl210)
.PROBE tran v(l1bl211)
.PROBE tran v(l1bl212)
.PROBE tran v(l1bl213)
.PROBE tran v(l1bl214)
.PROBE tran v(l1bl215)
.PROBE tran v(l1bl216)
.PROBE tran v(l1bl217)
.PROBE tran v(l1bl218)
.PROBE tran v(l1bl219)
.PROBE tran v(l1bl220)
.PROBE tran v(l1bl221)
.PROBE tran v(l1bl222)
.PROBE tran v(l1bl223)
.PROBE tran v(l1bl224)
.PROBE tran v(l1bl225)
.PROBE tran v(l1bl226)
.PROBE tran v(l1bl227)
.PROBE tran v(l1bl228)
.PROBE tran v(l1bl229)
.PROBE tran v(l1bl230)
.PROBE tran v(l1bl231)
.PROBE tran v(l1bl232)
.PROBE tran v(l1bl233)
.PROBE tran v(l1bl234)
.PROBE tran v(l1bl235)
.PROBE tran v(l1bl236)
.PROBE tran v(l1bl237)
.PROBE tran v(l1bl238)
.PROBE tran v(l1bl239)
.PROBE tran v(l1bl240)
.PROBE tran v(l1bl241)
.PROBE tran v(l1bl242)
.PROBE tran v(l1bl243)
.PROBE tran v(l1bl244)
.PROBE tran v(l1bl245)
.PROBE tran v(l1bl246)
.PROBE tran v(l1bl247)
.PROBE tran v(l1bl248)
.PROBE tran v(l1bl249)
.PROBE tran v(l1bl250)
.PROBE tran v(l1bl251)
.PROBE tran v(l1bl252)
.PROBE tran v(l1bl253)
.PROBE tran v(l1bl254)
.PROBE tran v(l1bl255)
.PROBE tran v(l1bl256)
.PROBE tran v(l1bl257)
.PROBE tran v(l1bl258)
.PROBE tran v(l1bl259)
.PROBE tran v(l1bl260)
.PROBE tran v(l1bl261)
.PROBE tran v(l1bl262)
.PROBE tran v(l1bl263)
.PROBE tran v(l1bl264)
.PROBE tran v(l1bl265)
.PROBE tran v(l1bl266)
.PROBE tran v(l1bl267)
.PROBE tran v(l1bl268)
.PROBE tran v(l1bl269)
.PROBE tran v(l1bl270)
.PROBE tran v(l1bl271)
.PROBE tran v(l1bl272)
.PROBE tran v(l1bl273)
.PROBE tran v(l1bl274)
.PROBE tran v(l1bl275)
.PROBE tran v(l1bl276)
.PROBE tran v(l1bl277)
.PROBE tran v(l1bl278)
.PROBE tran v(l1bl279)
.PROBE tran v(l1bl280)
.PROBE tran v(l1bl281)
.PROBE tran v(l1bl282)
.PROBE tran v(l1bl283)
.PROBE tran v(l1bl284)
.PROBE tran v(l1bl285)
.PROBE tran v(l1bl286)
.PROBE tran v(l1bl287)
.PROBE tran v(l1bl288)
.PROBE tran v(l1bl289)
.PROBE tran v(l1bl290)
.PROBE tran v(l1bl291)
.PROBE tran v(l1bl292)
.PROBE tran v(l1bl293)
.PROBE tran v(l1bl294)
.PROBE tran v(l1bl295)
.PROBE tran v(l1bl296)
.PROBE tran v(l1bl297)
.PROBE tran v(l1bl298)
.PROBE tran v(l1bl299)
.PROBE tran v(l1bl300)
.PROBE tran v(l1bl301)
.PROBE tran v(l1bl302)
.PROBE tran v(l1bl303)
.PROBE tran v(l1bl304)
.PROBE tran v(l1bl305)
.PROBE tran v(l1bl306)
.PROBE tran v(l1bl307)
.PROBE tran v(l1bl308)
.PROBE tran v(l1bl309)
.PROBE tran v(l1bl310)
.PROBE tran v(l1bl311)
.PROBE tran v(l1bl312)
.PROBE tran v(l1bl313)
.PROBE tran v(l1bl314)
.PROBE tran v(l1bl315)
.PROBE tran v(l1bl316)
.PROBE tran v(l1bl317)
.PROBE tran v(l1bl318)
.PROBE tran v(l1bl319)
.PROBE tran v(l1bl320)
.PROBE tran v(l1bl321)
.PROBE tran v(l1bl322)
.PROBE tran v(l1bl323)
.PROBE tran v(l1bl324)
.PROBE tran v(l1bl325)
.PROBE tran v(l1bl326)
.PROBE tran v(l1bl327)
.PROBE tran v(l1bl328)
.PROBE tran v(l1bl329)
.PROBE tran v(l1bl330)
.PROBE tran v(l1bl331)
.PROBE tran v(l1bl332)
.PROBE tran v(l1bl333)
.PROBE tran v(l1bl334)
.PROBE tran v(l1bl335)
.PROBE tran v(l1bl336)
.PROBE tran v(l1bl337)
.PROBE tran v(l1bl338)
.PROBE tran v(l1bl339)
.PROBE tran v(l1bl340)
.PROBE tran v(l1bl341)
.PROBE tran v(l1bl342)
.PROBE tran v(l1bl343)
.PROBE tran v(l1bl344)
.PROBE tran v(l1bl345)
.PROBE tran v(l1bl346)
.PROBE tran v(l1bl347)
.PROBE tran v(l1bl348)
.PROBE tran v(l1bl349)
.PROBE tran v(l1bl350)
.PROBE tran v(l1bl351)
.PROBE tran v(l1bl352)
.PROBE tran v(l1bl353)
.PROBE tran v(l1bl354)
.PROBE tran v(l1bl355)
.PROBE tran v(l1bl356)
.PROBE tran v(l1bl357)
.PROBE tran v(l1bl358)
.PROBE tran v(l1bl359)
.PROBE tran v(l1bl360)
.PROBE tran v(l1bl361)
.PROBE tran v(l1bl362)
.PROBE tran v(l1bl363)
.PROBE tran v(l1bl364)
.PROBE tran v(l1bl365)
.PROBE tran v(l1bl366)
.PROBE tran v(l1bl367)
.PROBE tran v(l1bl368)
.PROBE tran v(l1bl369)
.PROBE tran v(l1bl370)
.PROBE tran v(l1bl371)
.PROBE tran v(l1bl372)
.PROBE tran v(l1bl373)
.PROBE tran v(l1bl374)
.PROBE tran v(l1bl375)
.PROBE tran v(l1bl376)
.PROBE tran v(l1bl377)
.PROBE tran v(l1bl378)
.PROBE tran v(l1bl379)
.PROBE tran v(l1bl380)
.PROBE tran v(l1bl381)
.PROBE tran v(l1bl382)
.PROBE tran v(l1bl383)
.PROBE tran v(l1bl384)
.PROBE tran v(l1bl385)
.PROBE tran v(l1bl386)
.PROBE tran v(l1bl387)
.PROBE tran v(l1bl388)
.PROBE tran v(l1bl389)
.PROBE tran v(l1bl390)
.PROBE tran v(l1bl391)
.PROBE tran v(l1bl392)
.PROBE tran v(l1bl393)
.PROBE tran v(l1bl394)
.PROBE tran v(l1bl395)
.PROBE tran v(l1bl396)
.PROBE tran v(l1bl397)
.PROBE tran v(l1bl398)
.PROBE tran v(l1bl399)
.PROBE tran v(l1bl400)
.PROBE tran v(l1bl401)
.PROBE tran v(l1bl402)
.PROBE tran v(l1bl403)
.PROBE tran v(l1bl404)
.PROBE tran v(l1bl405)
.PROBE tran v(l1bl406)
.PROBE tran v(l1bl407)
.PROBE tran v(l1bl408)
.PROBE tran v(l1bl409)
.PROBE tran v(l1bl410)
.PROBE tran v(l1bl411)
.PROBE tran v(l1bl412)
.PROBE tran v(l1bl413)
.PROBE tran v(l1bl414)
.PROBE tran v(l1bl415)
.PROBE tran v(l1bl416)
.PROBE tran v(l1bl417)
.PROBE tran v(l1bl418)
.PROBE tran v(l1bl419)
.PROBE tran v(l1bl420)
.PROBE tran v(l1bl421)
.PROBE tran v(l1bl422)
.PROBE tran v(l1bl423)
.PROBE tran v(l1bl424)
.PROBE tran v(l1bl425)
.PROBE tran v(l1bl426)
.PROBE tran v(l1bl427)
.PROBE tran v(l1bl428)
.PROBE tran v(l1bl429)
.PROBE tran v(l1bl430)
.PROBE tran v(l1bl431)
.PROBE tran v(l1bl432)
.PROBE tran v(l1bl433)
.PROBE tran v(l1bl434)
.PROBE tran v(l1bl435)
.PROBE tran v(l1bl436)
.PROBE tran v(l1bl437)
.PROBE tran v(l1bl438)
.PROBE tran v(l1bl439)
.PROBE tran v(l1bl440)
.PROBE tran v(l1bl441)
.PROBE tran v(l1bl442)
.PROBE tran v(l1bl443)
.PROBE tran v(l1bl444)
.PROBE tran v(l1bl445)
.PROBE tran v(l1bl446)
.PROBE tran v(l1bl447)
.PROBE tran v(l1bl448)
.PROBE tran v(l1bl449)
.PROBE tran v(l1bl450)
.PROBE tran v(l1bl451)
.PROBE tran v(l1bl452)
.PROBE tran v(l1bl453)
.PROBE tran v(l1bl454)
.PROBE tran v(l1bl455)
.PROBE tran v(l1bl456)
.PROBE tran v(l1bl457)
.PROBE tran v(l1bl458)
.PROBE tran v(l1bl459)
.PROBE tran v(l1bl460)
.PROBE tran v(l1bl461)
.PROBE tran v(l1bl462)
.PROBE tran v(l1bl463)
.PROBE tran v(l1bl464)
.PROBE tran v(l1bl465)
.PROBE tran v(l1bl466)
.PROBE tran v(l1bl467)
.PROBE tran v(l1bl468)
.PROBE tran v(l1bl469)
.PROBE tran v(l1bl470)
.PROBE tran v(l1bl471)
.PROBE tran v(l1bl472)
.PROBE tran v(l1bl473)
.PROBE tran v(l1bl474)
.PROBE tran v(l1bl475)
.PROBE tran v(l1bl476)
.PROBE tran v(l1bl477)
.PROBE tran v(l1bl478)
.PROBE tran v(l1bl479)
.PROBE tran v(l1bl480)
.PROBE tran v(l1bl481)
.PROBE tran v(l1bl482)
.PROBE tran v(l1bl483)
.PROBE tran v(l1bl484)
.PROBE tran v(l1bl485)
.PROBE tran v(l1bl486)
.PROBE tran v(l1bl487)
.PROBE tran v(l1bl488)
.PROBE tran v(l1bl489)
.PROBE tran v(l1bl490)
.PROBE tran v(l1bl491)
.PROBE tran v(l1bl492)
.PROBE tran v(l1bl493)
.PROBE tran v(l1bl494)
.PROBE tran v(l1bl495)
.PROBE tran v(l1bl496)
.PROBE tran v(l1bl497)
.PROBE tran v(l1bl498)
.PROBE tran v(l1bl499)
.PROBE tran v(l1bl500)
.PROBE tran v(l1bl501)
.PROBE tran v(l1bl502)
.PROBE tran v(l1bl503)
.PROBE tran v(l1bl504)
.PROBE tran v(l1bl505)
.PROBE tran v(l1bl506)
.PROBE tran v(l1bl507)
.PROBE tran v(l1bl508)
.PROBE tran v(l1bl509)
.PROBE tran v(l1bl510)
.PROBE tran v(l1bl511)

.PROBE tran v(l2bl0)
.PROBE tran v(l2bl1)
.PROBE tran v(l2bl2)
.PROBE tran v(l2bl3)
.PROBE tran v(l2bl4)
.PROBE tran v(l2bl5)
.PROBE tran v(l2bl6)
.PROBE tran v(l2bl7)
.PROBE tran v(l2bl8)
.PROBE tran v(l2bl9)
.PROBE tran v(l2bl10)
.PROBE tran v(l2bl11)
.PROBE tran v(l2bl12)
.PROBE tran v(l2bl13)
.PROBE tran v(l2bl14)
.PROBE tran v(l2bl15)
.PROBE tran v(l2bl16)
.PROBE tran v(l2bl17)
.PROBE tran v(l2bl18)
.PROBE tran v(l2bl19)
.PROBE tran v(l2bl20)
.PROBE tran v(l2bl21)
.PROBE tran v(l2bl22)
.PROBE tran v(l2bl23)
.PROBE tran v(l2bl24)
.PROBE tran v(l2bl25)
.PROBE tran v(l2bl26)
.PROBE tran v(l2bl27)
.PROBE tran v(l2bl28)
.PROBE tran v(l2bl29)
.PROBE tran v(l2bl30)
.PROBE tran v(l2bl31)
.PROBE tran v(l2bl32)
.PROBE tran v(l2bl33)
.PROBE tran v(l2bl34)
.PROBE tran v(l2bl35)
.PROBE tran v(l2bl36)
.PROBE tran v(l2bl37)
.PROBE tran v(l2bl38)
.PROBE tran v(l2bl39)
.PROBE tran v(l2bl40)
.PROBE tran v(l2bl41)
.PROBE tran v(l2bl42)
.PROBE tran v(l2bl43)
.PROBE tran v(l2bl44)
.PROBE tran v(l2bl45)
.PROBE tran v(l2bl46)
.PROBE tran v(l2bl47)
.PROBE tran v(l2bl48)
.PROBE tran v(l2bl49)
.PROBE tran v(l2bl50)
.PROBE tran v(l2bl51)
.PROBE tran v(l2bl52)
.PROBE tran v(l2bl53)
.PROBE tran v(l2bl54)
.PROBE tran v(l2bl55)
.PROBE tran v(l2bl56)
.PROBE tran v(l2bl57)
.PROBE tran v(l2bl58)
.PROBE tran v(l2bl59)
.PROBE tran v(l2bl60)
.PROBE tran v(l2bl61)
.PROBE tran v(l2bl62)
.PROBE tran v(l2bl63)
.PROBE tran v(l2bl64)
.PROBE tran v(l2bl65)
.PROBE tran v(l2bl66)
.PROBE tran v(l2bl67)
.PROBE tran v(l2bl68)
.PROBE tran v(l2bl69)
.PROBE tran v(l2bl70)
.PROBE tran v(l2bl71)
.PROBE tran v(l2bl72)
.PROBE tran v(l2bl73)
.PROBE tran v(l2bl74)
.PROBE tran v(l2bl75)
.PROBE tran v(l2bl76)
.PROBE tran v(l2bl77)
.PROBE tran v(l2bl78)
.PROBE tran v(l2bl79)
.PROBE tran v(l2bl80)
.PROBE tran v(l2bl81)
.PROBE tran v(l2bl82)
.PROBE tran v(l2bl83)
.PROBE tran v(l2bl84)
.PROBE tran v(l2bl85)
.PROBE tran v(l2bl86)
.PROBE tran v(l2bl87)
.PROBE tran v(l2bl88)
.PROBE tran v(l2bl89)
.PROBE tran v(l2bl90)
.PROBE tran v(l2bl91)
.PROBE tran v(l2bl92)
.PROBE tran v(l2bl93)
.PROBE tran v(l2bl94)
.PROBE tran v(l2bl95)
.PROBE tran v(l2bl96)
.PROBE tran v(l2bl97)
.PROBE tran v(l2bl98)
.PROBE tran v(l2bl99)
.PROBE tran v(l2bl100)
.PROBE tran v(l2bl101)
.PROBE tran v(l2bl102)
.PROBE tran v(l2bl103)
.PROBE tran v(l2bl104)
.PROBE tran v(l2bl105)
.PROBE tran v(l2bl106)
.PROBE tran v(l2bl107)
.PROBE tran v(l2bl108)
.PROBE tran v(l2bl109)
.PROBE tran v(l2bl110)
.PROBE tran v(l2bl111)
.PROBE tran v(l2bl112)
.PROBE tran v(l2bl113)
.PROBE tran v(l2bl114)
.PROBE tran v(l2bl115)
.PROBE tran v(l2bl116)
.PROBE tran v(l2bl117)
.PROBE tran v(l2bl118)
.PROBE tran v(l2bl119)
.PROBE tran v(l2bl120)
.PROBE tran v(l2bl121)
.PROBE tran v(l2bl122)
.PROBE tran v(l2bl123)
.PROBE tran v(l2bl124)
.PROBE tran v(l2bl125)
.PROBE tran v(l2bl126)
.PROBE tran v(l2bl127)
.PROBE tran v(l2bl128)
.PROBE tran v(l2bl129)
.PROBE tran v(l2bl130)
.PROBE tran v(l2bl131)
.PROBE tran v(l2bl132)
.PROBE tran v(l2bl133)
.PROBE tran v(l2bl134)
.PROBE tran v(l2bl135)
.PROBE tran v(l2bl136)
.PROBE tran v(l2bl137)
.PROBE tran v(l2bl138)
.PROBE tran v(l2bl139)
.PROBE tran v(l2bl140)
.PROBE tran v(l2bl141)
.PROBE tran v(l2bl142)
.PROBE tran v(l2bl143)
.PROBE tran v(l2bl144)
.PROBE tran v(l2bl145)
.PROBE tran v(l2bl146)
.PROBE tran v(l2bl147)
.PROBE tran v(l2bl148)
.PROBE tran v(l2bl149)
.PROBE tran v(l2bl150)
.PROBE tran v(l2bl151)
.PROBE tran v(l2bl152)
.PROBE tran v(l2bl153)
.PROBE tran v(l2bl154)
.PROBE tran v(l2bl155)
.PROBE tran v(l2bl156)
.PROBE tran v(l2bl157)
.PROBE tran v(l2bl158)
.PROBE tran v(l2bl159)
.PROBE tran v(l2bl160)
.PROBE tran v(l2bl161)
.PROBE tran v(l2bl162)
.PROBE tran v(l2bl163)
.PROBE tran v(l2bl164)
.PROBE tran v(l2bl165)
.PROBE tran v(l2bl166)
.PROBE tran v(l2bl167)
.PROBE tran v(l2bl168)
.PROBE tran v(l2bl169)
.PROBE tran v(l2bl170)
.PROBE tran v(l2bl171)
.PROBE tran v(l2bl172)
.PROBE tran v(l2bl173)
.PROBE tran v(l2bl174)
.PROBE tran v(l2bl175)
.PROBE tran v(l2bl176)
.PROBE tran v(l2bl177)
.PROBE tran v(l2bl178)
.PROBE tran v(l2bl179)
.PROBE tran v(l2bl180)
.PROBE tran v(l2bl181)
.PROBE tran v(l2bl182)
.PROBE tran v(l2bl183)
.PROBE tran v(l2bl184)
.PROBE tran v(l2bl185)
.PROBE tran v(l2bl186)
.PROBE tran v(l2bl187)
.PROBE tran v(l2bl188)
.PROBE tran v(l2bl189)
.PROBE tran v(l2bl190)
.PROBE tran v(l2bl191)
.PROBE tran v(l2bl192)
.PROBE tran v(l2bl193)
.PROBE tran v(l2bl194)
.PROBE tran v(l2bl195)
.PROBE tran v(l2bl196)
.PROBE tran v(l2bl197)
.PROBE tran v(l2bl198)
.PROBE tran v(l2bl199)
.PROBE tran v(l2bl200)
.PROBE tran v(l2bl201)
.PROBE tran v(l2bl202)
.PROBE tran v(l2bl203)
.PROBE tran v(l2bl204)
.PROBE tran v(l2bl205)
.PROBE tran v(l2bl206)
.PROBE tran v(l2bl207)
.PROBE tran v(l2bl208)
.PROBE tran v(l2bl209)
.PROBE tran v(l2bl210)
.PROBE tran v(l2bl211)
.PROBE tran v(l2bl212)
.PROBE tran v(l2bl213)
.PROBE tran v(l2bl214)
.PROBE tran v(l2bl215)
.PROBE tran v(l2bl216)
.PROBE tran v(l2bl217)
.PROBE tran v(l2bl218)
.PROBE tran v(l2bl219)
.PROBE tran v(l2bl220)
.PROBE tran v(l2bl221)
.PROBE tran v(l2bl222)
.PROBE tran v(l2bl223)
.PROBE tran v(l2bl224)
.PROBE tran v(l2bl225)
.PROBE tran v(l2bl226)
.PROBE tran v(l2bl227)
.PROBE tran v(l2bl228)
.PROBE tran v(l2bl229)
.PROBE tran v(l2bl230)
.PROBE tran v(l2bl231)
.PROBE tran v(l2bl232)
.PROBE tran v(l2bl233)
.PROBE tran v(l2bl234)
.PROBE tran v(l2bl235)
.PROBE tran v(l2bl236)
.PROBE tran v(l2bl237)
.PROBE tran v(l2bl238)
.PROBE tran v(l2bl239)
.PROBE tran v(l2bl240)
.PROBE tran v(l2bl241)
.PROBE tran v(l2bl242)
.PROBE tran v(l2bl243)
.PROBE tran v(l2bl244)
.PROBE tran v(l2bl245)
.PROBE tran v(l2bl246)
.PROBE tran v(l2bl247)
.PROBE tran v(l2bl248)
.PROBE tran v(l2bl249)
.PROBE tran v(l2bl250)
.PROBE tran v(l2bl251)
.PROBE tran v(l2bl252)
.PROBE tran v(l2bl253)
.PROBE tran v(l2bl254)
.PROBE tran v(l2bl255)
.PROBE tran v(l2bl256)
.PROBE tran v(l2bl257)
.PROBE tran v(l2bl258)
.PROBE tran v(l2bl259)
.PROBE tran v(l2bl260)
.PROBE tran v(l2bl261)
.PROBE tran v(l2bl262)
.PROBE tran v(l2bl263)
.PROBE tran v(l2bl264)
.PROBE tran v(l2bl265)
.PROBE tran v(l2bl266)
.PROBE tran v(l2bl267)
.PROBE tran v(l2bl268)
.PROBE tran v(l2bl269)
.PROBE tran v(l2bl270)
.PROBE tran v(l2bl271)
.PROBE tran v(l2bl272)
.PROBE tran v(l2bl273)
.PROBE tran v(l2bl274)
.PROBE tran v(l2bl275)
.PROBE tran v(l2bl276)
.PROBE tran v(l2bl277)
.PROBE tran v(l2bl278)
.PROBE tran v(l2bl279)
.PROBE tran v(l2bl280)
.PROBE tran v(l2bl281)
.PROBE tran v(l2bl282)
.PROBE tran v(l2bl283)
.PROBE tran v(l2bl284)
.PROBE tran v(l2bl285)
.PROBE tran v(l2bl286)
.PROBE tran v(l2bl287)
.PROBE tran v(l2bl288)
.PROBE tran v(l2bl289)
.PROBE tran v(l2bl290)
.PROBE tran v(l2bl291)
.PROBE tran v(l2bl292)
.PROBE tran v(l2bl293)
.PROBE tran v(l2bl294)
.PROBE tran v(l2bl295)
.PROBE tran v(l2bl296)
.PROBE tran v(l2bl297)
.PROBE tran v(l2bl298)
.PROBE tran v(l2bl299)
.PROBE tran v(l2bl300)
.PROBE tran v(l2bl301)
.PROBE tran v(l2bl302)
.PROBE tran v(l2bl303)
.PROBE tran v(l2bl304)
.PROBE tran v(l2bl305)
.PROBE tran v(l2bl306)
.PROBE tran v(l2bl307)
.PROBE tran v(l2bl308)
.PROBE tran v(l2bl309)
.PROBE tran v(l2bl310)
.PROBE tran v(l2bl311)
.PROBE tran v(l2bl312)
.PROBE tran v(l2bl313)
.PROBE tran v(l2bl314)
.PROBE tran v(l2bl315)
.PROBE tran v(l2bl316)
.PROBE tran v(l2bl317)
.PROBE tran v(l2bl318)
.PROBE tran v(l2bl319)
.PROBE tran v(l2bl320)
.PROBE tran v(l2bl321)
.PROBE tran v(l2bl322)
.PROBE tran v(l2bl323)
.PROBE tran v(l2bl324)
.PROBE tran v(l2bl325)
.PROBE tran v(l2bl326)
.PROBE tran v(l2bl327)
.PROBE tran v(l2bl328)
.PROBE tran v(l2bl329)
.PROBE tran v(l2bl330)
.PROBE tran v(l2bl331)
.PROBE tran v(l2bl332)
.PROBE tran v(l2bl333)
.PROBE tran v(l2bl334)
.PROBE tran v(l2bl335)
.PROBE tran v(l2bl336)
.PROBE tran v(l2bl337)
.PROBE tran v(l2bl338)
.PROBE tran v(l2bl339)
.PROBE tran v(l2bl340)
.PROBE tran v(l2bl341)
.PROBE tran v(l2bl342)
.PROBE tran v(l2bl343)
.PROBE tran v(l2bl344)
.PROBE tran v(l2bl345)
.PROBE tran v(l2bl346)
.PROBE tran v(l2bl347)
.PROBE tran v(l2bl348)
.PROBE tran v(l2bl349)
.PROBE tran v(l2bl350)
.PROBE tran v(l2bl351)
.PROBE tran v(l2bl352)
.PROBE tran v(l2bl353)
.PROBE tran v(l2bl354)
.PROBE tran v(l2bl355)
.PROBE tran v(l2bl356)
.PROBE tran v(l2bl357)
.PROBE tran v(l2bl358)
.PROBE tran v(l2bl359)
.PROBE tran v(l2bl360)
.PROBE tran v(l2bl361)
.PROBE tran v(l2bl362)
.PROBE tran v(l2bl363)
.PROBE tran v(l2bl364)
.PROBE tran v(l2bl365)
.PROBE tran v(l2bl366)
.PROBE tran v(l2bl367)
.PROBE tran v(l2bl368)
.PROBE tran v(l2bl369)
.PROBE tran v(l2bl370)
.PROBE tran v(l2bl371)
.PROBE tran v(l2bl372)
.PROBE tran v(l2bl373)
.PROBE tran v(l2bl374)
.PROBE tran v(l2bl375)
.PROBE tran v(l2bl376)
.PROBE tran v(l2bl377)
.PROBE tran v(l2bl378)
.PROBE tran v(l2bl379)
.PROBE tran v(l2bl380)
.PROBE tran v(l2bl381)
.PROBE tran v(l2bl382)
.PROBE tran v(l2bl383)
.PROBE tran v(l2bl384)
.PROBE tran v(l2bl385)
.PROBE tran v(l2bl386)
.PROBE tran v(l2bl387)
.PROBE tran v(l2bl388)
.PROBE tran v(l2bl389)
.PROBE tran v(l2bl390)
.PROBE tran v(l2bl391)
.PROBE tran v(l2bl392)
.PROBE tran v(l2bl393)
.PROBE tran v(l2bl394)
.PROBE tran v(l2bl395)
.PROBE tran v(l2bl396)
.PROBE tran v(l2bl397)
.PROBE tran v(l2bl398)
.PROBE tran v(l2bl399)
.PROBE tran v(l2bl400)
.PROBE tran v(l2bl401)
.PROBE tran v(l2bl402)
.PROBE tran v(l2bl403)
.PROBE tran v(l2bl404)
.PROBE tran v(l2bl405)
.PROBE tran v(l2bl406)
.PROBE tran v(l2bl407)
.PROBE tran v(l2bl408)
.PROBE tran v(l2bl409)
.PROBE tran v(l2bl410)
.PROBE tran v(l2bl411)
.PROBE tran v(l2bl412)
.PROBE tran v(l2bl413)
.PROBE tran v(l2bl414)
.PROBE tran v(l2bl415)
.PROBE tran v(l2bl416)
.PROBE tran v(l2bl417)
.PROBE tran v(l2bl418)
.PROBE tran v(l2bl419)
.PROBE tran v(l2bl420)
.PROBE tran v(l2bl421)
.PROBE tran v(l2bl422)
.PROBE tran v(l2bl423)
.PROBE tran v(l2bl424)
.PROBE tran v(l2bl425)
.PROBE tran v(l2bl426)
.PROBE tran v(l2bl427)
.PROBE tran v(l2bl428)
.PROBE tran v(l2bl429)
.PROBE tran v(l2bl430)
.PROBE tran v(l2bl431)
.PROBE tran v(l2bl432)
.PROBE tran v(l2bl433)
.PROBE tran v(l2bl434)
.PROBE tran v(l2bl435)
.PROBE tran v(l2bl436)
.PROBE tran v(l2bl437)
.PROBE tran v(l2bl438)
.PROBE tran v(l2bl439)
.PROBE tran v(l2bl440)
.PROBE tran v(l2bl441)
.PROBE tran v(l2bl442)
.PROBE tran v(l2bl443)
.PROBE tran v(l2bl444)
.PROBE tran v(l2bl445)
.PROBE tran v(l2bl446)
.PROBE tran v(l2bl447)
.PROBE tran v(l2bl448)
.PROBE tran v(l2bl449)
.PROBE tran v(l2bl450)
.PROBE tran v(l2bl451)
.PROBE tran v(l2bl452)
.PROBE tran v(l2bl453)
.PROBE tran v(l2bl454)
.PROBE tran v(l2bl455)
.PROBE tran v(l2bl456)
.PROBE tran v(l2bl457)
.PROBE tran v(l2bl458)
.PROBE tran v(l2bl459)
.PROBE tran v(l2bl460)
.PROBE tran v(l2bl461)
.PROBE tran v(l2bl462)
.PROBE tran v(l2bl463)
.PROBE tran v(l2bl464)
.PROBE tran v(l2bl465)
.PROBE tran v(l2bl466)
.PROBE tran v(l2bl467)
.PROBE tran v(l2bl468)
.PROBE tran v(l2bl469)
.PROBE tran v(l2bl470)
.PROBE tran v(l2bl471)
.PROBE tran v(l2bl472)
.PROBE tran v(l2bl473)
.PROBE tran v(l2bl474)
.PROBE tran v(l2bl475)
.PROBE tran v(l2bl476)
.PROBE tran v(l2bl477)
.PROBE tran v(l2bl478)
.PROBE tran v(l2bl479)
.PROBE tran v(l2bl480)
.PROBE tran v(l2bl481)
.PROBE tran v(l2bl482)
.PROBE tran v(l2bl483)
.PROBE tran v(l2bl484)
.PROBE tran v(l2bl485)
.PROBE tran v(l2bl486)
.PROBE tran v(l2bl487)
.PROBE tran v(l2bl488)
.PROBE tran v(l2bl489)
.PROBE tran v(l2bl490)
.PROBE tran v(l2bl491)
.PROBE tran v(l2bl492)
.PROBE tran v(l2bl493)
.PROBE tran v(l2bl494)
.PROBE tran v(l2bl495)
.PROBE tran v(l2bl496)
.PROBE tran v(l2bl497)
.PROBE tran v(l2bl498)
.PROBE tran v(l2bl499)
.PROBE tran v(l2bl500)
.PROBE tran v(l2bl501)
.PROBE tran v(l2bl502)
.PROBE tran v(l2bl503)
.PROBE tran v(l2bl504)
.PROBE tran v(l2bl505)
.PROBE tran v(l2bl506)
.PROBE tran v(l2bl507)
.PROBE tran v(l2bl508)
.PROBE tran v(l2bl509)
.PROBE tran v(l2bl510)
.PROBE tran v(l2bl511)

.measure tran avgvall0bl0 AVG v(l0bl0) FROM = 0ns TO =1ns
.measure tran avgvall0bl1 AVG v(l0bl1) FROM = 0ns TO =1ns
.measure tran avgvall0bl2 AVG v(l0bl2) FROM = 0ns TO =1ns
.measure tran avgvall0bl3 AVG v(l0bl3) FROM = 0ns TO =1ns
.measure tran avgvall0bl4 AVG v(l0bl4) FROM = 0ns TO =1ns
.measure tran avgvall0bl5 AVG v(l0bl5) FROM = 0ns TO =1ns
.measure tran avgvall0bl6 AVG v(l0bl6) FROM = 0ns TO =1ns
.measure tran avgvall0bl7 AVG v(l0bl7) FROM = 0ns TO =1ns
.measure tran avgvall0bl8 AVG v(l0bl8) FROM = 0ns TO =1ns
.measure tran avgvall0bl9 AVG v(l0bl9) FROM = 0ns TO =1ns
.measure tran avgvall0bl10 AVG v(l0bl10) FROM = 0ns TO =1ns
.measure tran avgvall0bl11 AVG v(l0bl11) FROM = 0ns TO =1ns
.measure tran avgvall0bl12 AVG v(l0bl12) FROM = 0ns TO =1ns
.measure tran avgvall0bl13 AVG v(l0bl13) FROM = 0ns TO =1ns
.measure tran avgvall0bl14 AVG v(l0bl14) FROM = 0ns TO =1ns
.measure tran avgvall0bl15 AVG v(l0bl15) FROM = 0ns TO =1ns
.measure tran avgvall0bl16 AVG v(l0bl16) FROM = 0ns TO =1ns
.measure tran avgvall0bl17 AVG v(l0bl17) FROM = 0ns TO =1ns
.measure tran avgvall0bl18 AVG v(l0bl18) FROM = 0ns TO =1ns
.measure tran avgvall0bl19 AVG v(l0bl19) FROM = 0ns TO =1ns
.measure tran avgvall0bl20 AVG v(l0bl20) FROM = 0ns TO =1ns
.measure tran avgvall0bl21 AVG v(l0bl21) FROM = 0ns TO =1ns
.measure tran avgvall0bl22 AVG v(l0bl22) FROM = 0ns TO =1ns
.measure tran avgvall0bl23 AVG v(l0bl23) FROM = 0ns TO =1ns
.measure tran avgvall0bl24 AVG v(l0bl24) FROM = 0ns TO =1ns
.measure tran avgvall0bl25 AVG v(l0bl25) FROM = 0ns TO =1ns
.measure tran avgvall0bl26 AVG v(l0bl26) FROM = 0ns TO =1ns
.measure tran avgvall0bl27 AVG v(l0bl27) FROM = 0ns TO =1ns
.measure tran avgvall0bl28 AVG v(l0bl28) FROM = 0ns TO =1ns
.measure tran avgvall0bl29 AVG v(l0bl29) FROM = 0ns TO =1ns
.measure tran avgvall0bl30 AVG v(l0bl30) FROM = 0ns TO =1ns
.measure tran avgvall0bl31 AVG v(l0bl31) FROM = 0ns TO =1ns
.measure tran avgvall0bl32 AVG v(l0bl32) FROM = 0ns TO =1ns
.measure tran avgvall0bl33 AVG v(l0bl33) FROM = 0ns TO =1ns
.measure tran avgvall0bl34 AVG v(l0bl34) FROM = 0ns TO =1ns
.measure tran avgvall0bl35 AVG v(l0bl35) FROM = 0ns TO =1ns
.measure tran avgvall0bl36 AVG v(l0bl36) FROM = 0ns TO =1ns
.measure tran avgvall0bl37 AVG v(l0bl37) FROM = 0ns TO =1ns
.measure tran avgvall0bl38 AVG v(l0bl38) FROM = 0ns TO =1ns
.measure tran avgvall0bl39 AVG v(l0bl39) FROM = 0ns TO =1ns
.measure tran avgvall0bl40 AVG v(l0bl40) FROM = 0ns TO =1ns
.measure tran avgvall0bl41 AVG v(l0bl41) FROM = 0ns TO =1ns
.measure tran avgvall0bl42 AVG v(l0bl42) FROM = 0ns TO =1ns
.measure tran avgvall0bl43 AVG v(l0bl43) FROM = 0ns TO =1ns
.measure tran avgvall0bl44 AVG v(l0bl44) FROM = 0ns TO =1ns
.measure tran avgvall0bl45 AVG v(l0bl45) FROM = 0ns TO =1ns
.measure tran avgvall0bl46 AVG v(l0bl46) FROM = 0ns TO =1ns
.measure tran avgvall0bl47 AVG v(l0bl47) FROM = 0ns TO =1ns
.measure tran avgvall0bl48 AVG v(l0bl48) FROM = 0ns TO =1ns
.measure tran avgvall0bl49 AVG v(l0bl49) FROM = 0ns TO =1ns
.measure tran avgvall0bl50 AVG v(l0bl50) FROM = 0ns TO =1ns
.measure tran avgvall0bl51 AVG v(l0bl51) FROM = 0ns TO =1ns
.measure tran avgvall0bl52 AVG v(l0bl52) FROM = 0ns TO =1ns
.measure tran avgvall0bl53 AVG v(l0bl53) FROM = 0ns TO =1ns
.measure tran avgvall0bl54 AVG v(l0bl54) FROM = 0ns TO =1ns
.measure tran avgvall0bl55 AVG v(l0bl55) FROM = 0ns TO =1ns
.measure tran avgvall0bl56 AVG v(l0bl56) FROM = 0ns TO =1ns
.measure tran avgvall0bl57 AVG v(l0bl57) FROM = 0ns TO =1ns
.measure tran avgvall0bl58 AVG v(l0bl58) FROM = 0ns TO =1ns
.measure tran avgvall0bl59 AVG v(l0bl59) FROM = 0ns TO =1ns
.measure tran avgvall0bl60 AVG v(l0bl60) FROM = 0ns TO =1ns
.measure tran avgvall0bl61 AVG v(l0bl61) FROM = 0ns TO =1ns
.measure tran avgvall0bl62 AVG v(l0bl62) FROM = 0ns TO =1ns
.measure tran avgvall0bl63 AVG v(l0bl63) FROM = 0ns TO =1ns
.measure tran avgvall0bl64 AVG v(l0bl64) FROM = 0ns TO =1ns
.measure tran avgvall0bl65 AVG v(l0bl65) FROM = 0ns TO =1ns
.measure tran avgvall0bl66 AVG v(l0bl66) FROM = 0ns TO =1ns
.measure tran avgvall0bl67 AVG v(l0bl67) FROM = 0ns TO =1ns
.measure tran avgvall0bl68 AVG v(l0bl68) FROM = 0ns TO =1ns
.measure tran avgvall0bl69 AVG v(l0bl69) FROM = 0ns TO =1ns
.measure tran avgvall0bl70 AVG v(l0bl70) FROM = 0ns TO =1ns
.measure tran avgvall0bl71 AVG v(l0bl71) FROM = 0ns TO =1ns
.measure tran avgvall0bl72 AVG v(l0bl72) FROM = 0ns TO =1ns
.measure tran avgvall0bl73 AVG v(l0bl73) FROM = 0ns TO =1ns
.measure tran avgvall0bl74 AVG v(l0bl74) FROM = 0ns TO =1ns
.measure tran avgvall0bl75 AVG v(l0bl75) FROM = 0ns TO =1ns
.measure tran avgvall0bl76 AVG v(l0bl76) FROM = 0ns TO =1ns
.measure tran avgvall0bl77 AVG v(l0bl77) FROM = 0ns TO =1ns
.measure tran avgvall0bl78 AVG v(l0bl78) FROM = 0ns TO =1ns
.measure tran avgvall0bl79 AVG v(l0bl79) FROM = 0ns TO =1ns
.measure tran avgvall0bl80 AVG v(l0bl80) FROM = 0ns TO =1ns
.measure tran avgvall0bl81 AVG v(l0bl81) FROM = 0ns TO =1ns
.measure tran avgvall0bl82 AVG v(l0bl82) FROM = 0ns TO =1ns
.measure tran avgvall0bl83 AVG v(l0bl83) FROM = 0ns TO =1ns
.measure tran avgvall0bl84 AVG v(l0bl84) FROM = 0ns TO =1ns
.measure tran avgvall0bl85 AVG v(l0bl85) FROM = 0ns TO =1ns
.measure tran avgvall0bl86 AVG v(l0bl86) FROM = 0ns TO =1ns
.measure tran avgvall0bl87 AVG v(l0bl87) FROM = 0ns TO =1ns
.measure tran avgvall0bl88 AVG v(l0bl88) FROM = 0ns TO =1ns
.measure tran avgvall0bl89 AVG v(l0bl89) FROM = 0ns TO =1ns
.measure tran avgvall0bl90 AVG v(l0bl90) FROM = 0ns TO =1ns
.measure tran avgvall0bl91 AVG v(l0bl91) FROM = 0ns TO =1ns
.measure tran avgvall0bl92 AVG v(l0bl92) FROM = 0ns TO =1ns
.measure tran avgvall0bl93 AVG v(l0bl93) FROM = 0ns TO =1ns
.measure tran avgvall0bl94 AVG v(l0bl94) FROM = 0ns TO =1ns
.measure tran avgvall0bl95 AVG v(l0bl95) FROM = 0ns TO =1ns
.measure tran avgvall0bl96 AVG v(l0bl96) FROM = 0ns TO =1ns
.measure tran avgvall0bl97 AVG v(l0bl97) FROM = 0ns TO =1ns
.measure tran avgvall0bl98 AVG v(l0bl98) FROM = 0ns TO =1ns
.measure tran avgvall0bl99 AVG v(l0bl99) FROM = 0ns TO =1ns
.measure tran avgvall0bl100 AVG v(l0bl100) FROM = 0ns TO =1ns
.measure tran avgvall0bl101 AVG v(l0bl101) FROM = 0ns TO =1ns
.measure tran avgvall0bl102 AVG v(l0bl102) FROM = 0ns TO =1ns
.measure tran avgvall0bl103 AVG v(l0bl103) FROM = 0ns TO =1ns
.measure tran avgvall0bl104 AVG v(l0bl104) FROM = 0ns TO =1ns
.measure tran avgvall0bl105 AVG v(l0bl105) FROM = 0ns TO =1ns
.measure tran avgvall0bl106 AVG v(l0bl106) FROM = 0ns TO =1ns
.measure tran avgvall0bl107 AVG v(l0bl107) FROM = 0ns TO =1ns
.measure tran avgvall0bl108 AVG v(l0bl108) FROM = 0ns TO =1ns
.measure tran avgvall0bl109 AVG v(l0bl109) FROM = 0ns TO =1ns
.measure tran avgvall0bl110 AVG v(l0bl110) FROM = 0ns TO =1ns
.measure tran avgvall0bl111 AVG v(l0bl111) FROM = 0ns TO =1ns
.measure tran avgvall0bl112 AVG v(l0bl112) FROM = 0ns TO =1ns
.measure tran avgvall0bl113 AVG v(l0bl113) FROM = 0ns TO =1ns
.measure tran avgvall0bl114 AVG v(l0bl114) FROM = 0ns TO =1ns
.measure tran avgvall0bl115 AVG v(l0bl115) FROM = 0ns TO =1ns
.measure tran avgvall0bl116 AVG v(l0bl116) FROM = 0ns TO =1ns
.measure tran avgvall0bl117 AVG v(l0bl117) FROM = 0ns TO =1ns
.measure tran avgvall0bl118 AVG v(l0bl118) FROM = 0ns TO =1ns
.measure tran avgvall0bl119 AVG v(l0bl119) FROM = 0ns TO =1ns
.measure tran avgvall0bl120 AVG v(l0bl120) FROM = 0ns TO =1ns
.measure tran avgvall0bl121 AVG v(l0bl121) FROM = 0ns TO =1ns
.measure tran avgvall0bl122 AVG v(l0bl122) FROM = 0ns TO =1ns
.measure tran avgvall0bl123 AVG v(l0bl123) FROM = 0ns TO =1ns
.measure tran avgvall0bl124 AVG v(l0bl124) FROM = 0ns TO =1ns
.measure tran avgvall0bl125 AVG v(l0bl125) FROM = 0ns TO =1ns
.measure tran avgvall0bl126 AVG v(l0bl126) FROM = 0ns TO =1ns
.measure tran avgvall0bl127 AVG v(l0bl127) FROM = 0ns TO =1ns
.measure tran avgvall0bl128 AVG v(l0bl128) FROM = 0ns TO =1ns
.measure tran avgvall0bl129 AVG v(l0bl129) FROM = 0ns TO =1ns
.measure tran avgvall0bl130 AVG v(l0bl130) FROM = 0ns TO =1ns
.measure tran avgvall0bl131 AVG v(l0bl131) FROM = 0ns TO =1ns
.measure tran avgvall0bl132 AVG v(l0bl132) FROM = 0ns TO =1ns
.measure tran avgvall0bl133 AVG v(l0bl133) FROM = 0ns TO =1ns
.measure tran avgvall0bl134 AVG v(l0bl134) FROM = 0ns TO =1ns
.measure tran avgvall0bl135 AVG v(l0bl135) FROM = 0ns TO =1ns
.measure tran avgvall0bl136 AVG v(l0bl136) FROM = 0ns TO =1ns
.measure tran avgvall0bl137 AVG v(l0bl137) FROM = 0ns TO =1ns
.measure tran avgvall0bl138 AVG v(l0bl138) FROM = 0ns TO =1ns
.measure tran avgvall0bl139 AVG v(l0bl139) FROM = 0ns TO =1ns
.measure tran avgvall0bl140 AVG v(l0bl140) FROM = 0ns TO =1ns
.measure tran avgvall0bl141 AVG v(l0bl141) FROM = 0ns TO =1ns
.measure tran avgvall0bl142 AVG v(l0bl142) FROM = 0ns TO =1ns
.measure tran avgvall0bl143 AVG v(l0bl143) FROM = 0ns TO =1ns
.measure tran avgvall0bl144 AVG v(l0bl144) FROM = 0ns TO =1ns
.measure tran avgvall0bl145 AVG v(l0bl145) FROM = 0ns TO =1ns
.measure tran avgvall0bl146 AVG v(l0bl146) FROM = 0ns TO =1ns
.measure tran avgvall0bl147 AVG v(l0bl147) FROM = 0ns TO =1ns
.measure tran avgvall0bl148 AVG v(l0bl148) FROM = 0ns TO =1ns
.measure tran avgvall0bl149 AVG v(l0bl149) FROM = 0ns TO =1ns
.measure tran avgvall0bl150 AVG v(l0bl150) FROM = 0ns TO =1ns
.measure tran avgvall0bl151 AVG v(l0bl151) FROM = 0ns TO =1ns
.measure tran avgvall0bl152 AVG v(l0bl152) FROM = 0ns TO =1ns
.measure tran avgvall0bl153 AVG v(l0bl153) FROM = 0ns TO =1ns
.measure tran avgvall0bl154 AVG v(l0bl154) FROM = 0ns TO =1ns
.measure tran avgvall0bl155 AVG v(l0bl155) FROM = 0ns TO =1ns
.measure tran avgvall0bl156 AVG v(l0bl156) FROM = 0ns TO =1ns
.measure tran avgvall0bl157 AVG v(l0bl157) FROM = 0ns TO =1ns
.measure tran avgvall0bl158 AVG v(l0bl158) FROM = 0ns TO =1ns
.measure tran avgvall0bl159 AVG v(l0bl159) FROM = 0ns TO =1ns
.measure tran avgvall0bl160 AVG v(l0bl160) FROM = 0ns TO =1ns
.measure tran avgvall0bl161 AVG v(l0bl161) FROM = 0ns TO =1ns
.measure tran avgvall0bl162 AVG v(l0bl162) FROM = 0ns TO =1ns
.measure tran avgvall0bl163 AVG v(l0bl163) FROM = 0ns TO =1ns
.measure tran avgvall0bl164 AVG v(l0bl164) FROM = 0ns TO =1ns
.measure tran avgvall0bl165 AVG v(l0bl165) FROM = 0ns TO =1ns
.measure tran avgvall0bl166 AVG v(l0bl166) FROM = 0ns TO =1ns
.measure tran avgvall0bl167 AVG v(l0bl167) FROM = 0ns TO =1ns
.measure tran avgvall0bl168 AVG v(l0bl168) FROM = 0ns TO =1ns
.measure tran avgvall0bl169 AVG v(l0bl169) FROM = 0ns TO =1ns
.measure tran avgvall0bl170 AVG v(l0bl170) FROM = 0ns TO =1ns
.measure tran avgvall0bl171 AVG v(l0bl171) FROM = 0ns TO =1ns
.measure tran avgvall0bl172 AVG v(l0bl172) FROM = 0ns TO =1ns
.measure tran avgvall0bl173 AVG v(l0bl173) FROM = 0ns TO =1ns
.measure tran avgvall0bl174 AVG v(l0bl174) FROM = 0ns TO =1ns
.measure tran avgvall0bl175 AVG v(l0bl175) FROM = 0ns TO =1ns
.measure tran avgvall0bl176 AVG v(l0bl176) FROM = 0ns TO =1ns
.measure tran avgvall0bl177 AVG v(l0bl177) FROM = 0ns TO =1ns
.measure tran avgvall0bl178 AVG v(l0bl178) FROM = 0ns TO =1ns
.measure tran avgvall0bl179 AVG v(l0bl179) FROM = 0ns TO =1ns
.measure tran avgvall0bl180 AVG v(l0bl180) FROM = 0ns TO =1ns
.measure tran avgvall0bl181 AVG v(l0bl181) FROM = 0ns TO =1ns
.measure tran avgvall0bl182 AVG v(l0bl182) FROM = 0ns TO =1ns
.measure tran avgvall0bl183 AVG v(l0bl183) FROM = 0ns TO =1ns
.measure tran avgvall0bl184 AVG v(l0bl184) FROM = 0ns TO =1ns
.measure tran avgvall0bl185 AVG v(l0bl185) FROM = 0ns TO =1ns
.measure tran avgvall0bl186 AVG v(l0bl186) FROM = 0ns TO =1ns
.measure tran avgvall0bl187 AVG v(l0bl187) FROM = 0ns TO =1ns
.measure tran avgvall0bl188 AVG v(l0bl188) FROM = 0ns TO =1ns
.measure tran avgvall0bl189 AVG v(l0bl189) FROM = 0ns TO =1ns
.measure tran avgvall0bl190 AVG v(l0bl190) FROM = 0ns TO =1ns
.measure tran avgvall0bl191 AVG v(l0bl191) FROM = 0ns TO =1ns
.measure tran avgvall0bl192 AVG v(l0bl192) FROM = 0ns TO =1ns
.measure tran avgvall0bl193 AVG v(l0bl193) FROM = 0ns TO =1ns
.measure tran avgvall0bl194 AVG v(l0bl194) FROM = 0ns TO =1ns
.measure tran avgvall0bl195 AVG v(l0bl195) FROM = 0ns TO =1ns
.measure tran avgvall0bl196 AVG v(l0bl196) FROM = 0ns TO =1ns
.measure tran avgvall0bl197 AVG v(l0bl197) FROM = 0ns TO =1ns
.measure tran avgvall0bl198 AVG v(l0bl198) FROM = 0ns TO =1ns
.measure tran avgvall0bl199 AVG v(l0bl199) FROM = 0ns TO =1ns
.measure tran avgvall0bl200 AVG v(l0bl200) FROM = 0ns TO =1ns
.measure tran avgvall0bl201 AVG v(l0bl201) FROM = 0ns TO =1ns
.measure tran avgvall0bl202 AVG v(l0bl202) FROM = 0ns TO =1ns
.measure tran avgvall0bl203 AVG v(l0bl203) FROM = 0ns TO =1ns
.measure tran avgvall0bl204 AVG v(l0bl204) FROM = 0ns TO =1ns
.measure tran avgvall0bl205 AVG v(l0bl205) FROM = 0ns TO =1ns
.measure tran avgvall0bl206 AVG v(l0bl206) FROM = 0ns TO =1ns
.measure tran avgvall0bl207 AVG v(l0bl207) FROM = 0ns TO =1ns
.measure tran avgvall0bl208 AVG v(l0bl208) FROM = 0ns TO =1ns
.measure tran avgvall0bl209 AVG v(l0bl209) FROM = 0ns TO =1ns
.measure tran avgvall0bl210 AVG v(l0bl210) FROM = 0ns TO =1ns
.measure tran avgvall0bl211 AVG v(l0bl211) FROM = 0ns TO =1ns
.measure tran avgvall0bl212 AVG v(l0bl212) FROM = 0ns TO =1ns
.measure tran avgvall0bl213 AVG v(l0bl213) FROM = 0ns TO =1ns
.measure tran avgvall0bl214 AVG v(l0bl214) FROM = 0ns TO =1ns
.measure tran avgvall0bl215 AVG v(l0bl215) FROM = 0ns TO =1ns
.measure tran avgvall0bl216 AVG v(l0bl216) FROM = 0ns TO =1ns
.measure tran avgvall0bl217 AVG v(l0bl217) FROM = 0ns TO =1ns
.measure tran avgvall0bl218 AVG v(l0bl218) FROM = 0ns TO =1ns
.measure tran avgvall0bl219 AVG v(l0bl219) FROM = 0ns TO =1ns
.measure tran avgvall0bl220 AVG v(l0bl220) FROM = 0ns TO =1ns
.measure tran avgvall0bl221 AVG v(l0bl221) FROM = 0ns TO =1ns
.measure tran avgvall0bl222 AVG v(l0bl222) FROM = 0ns TO =1ns
.measure tran avgvall0bl223 AVG v(l0bl223) FROM = 0ns TO =1ns
.measure tran avgvall0bl224 AVG v(l0bl224) FROM = 0ns TO =1ns
.measure tran avgvall0bl225 AVG v(l0bl225) FROM = 0ns TO =1ns
.measure tran avgvall0bl226 AVG v(l0bl226) FROM = 0ns TO =1ns
.measure tran avgvall0bl227 AVG v(l0bl227) FROM = 0ns TO =1ns
.measure tran avgvall0bl228 AVG v(l0bl228) FROM = 0ns TO =1ns
.measure tran avgvall0bl229 AVG v(l0bl229) FROM = 0ns TO =1ns
.measure tran avgvall0bl230 AVG v(l0bl230) FROM = 0ns TO =1ns
.measure tran avgvall0bl231 AVG v(l0bl231) FROM = 0ns TO =1ns
.measure tran avgvall0bl232 AVG v(l0bl232) FROM = 0ns TO =1ns
.measure tran avgvall0bl233 AVG v(l0bl233) FROM = 0ns TO =1ns
.measure tran avgvall0bl234 AVG v(l0bl234) FROM = 0ns TO =1ns
.measure tran avgvall0bl235 AVG v(l0bl235) FROM = 0ns TO =1ns
.measure tran avgvall0bl236 AVG v(l0bl236) FROM = 0ns TO =1ns
.measure tran avgvall0bl237 AVG v(l0bl237) FROM = 0ns TO =1ns
.measure tran avgvall0bl238 AVG v(l0bl238) FROM = 0ns TO =1ns
.measure tran avgvall0bl239 AVG v(l0bl239) FROM = 0ns TO =1ns
.measure tran avgvall0bl240 AVG v(l0bl240) FROM = 0ns TO =1ns
.measure tran avgvall0bl241 AVG v(l0bl241) FROM = 0ns TO =1ns
.measure tran avgvall0bl242 AVG v(l0bl242) FROM = 0ns TO =1ns
.measure tran avgvall0bl243 AVG v(l0bl243) FROM = 0ns TO =1ns
.measure tran avgvall0bl244 AVG v(l0bl244) FROM = 0ns TO =1ns
.measure tran avgvall0bl245 AVG v(l0bl245) FROM = 0ns TO =1ns
.measure tran avgvall0bl246 AVG v(l0bl246) FROM = 0ns TO =1ns
.measure tran avgvall0bl247 AVG v(l0bl247) FROM = 0ns TO =1ns
.measure tran avgvall0bl248 AVG v(l0bl248) FROM = 0ns TO =1ns
.measure tran avgvall0bl249 AVG v(l0bl249) FROM = 0ns TO =1ns
.measure tran avgvall0bl250 AVG v(l0bl250) FROM = 0ns TO =1ns
.measure tran avgvall0bl251 AVG v(l0bl251) FROM = 0ns TO =1ns
.measure tran avgvall0bl252 AVG v(l0bl252) FROM = 0ns TO =1ns
.measure tran avgvall0bl253 AVG v(l0bl253) FROM = 0ns TO =1ns
.measure tran avgvall0bl254 AVG v(l0bl254) FROM = 0ns TO =1ns
.measure tran avgvall0bl255 AVG v(l0bl255) FROM = 0ns TO =1ns
.measure tran avgvall0bl256 AVG v(l0bl256) FROM = 0ns TO =1ns
.measure tran avgvall0bl257 AVG v(l0bl257) FROM = 0ns TO =1ns
.measure tran avgvall0bl258 AVG v(l0bl258) FROM = 0ns TO =1ns
.measure tran avgvall0bl259 AVG v(l0bl259) FROM = 0ns TO =1ns
.measure tran avgvall0bl260 AVG v(l0bl260) FROM = 0ns TO =1ns
.measure tran avgvall0bl261 AVG v(l0bl261) FROM = 0ns TO =1ns
.measure tran avgvall0bl262 AVG v(l0bl262) FROM = 0ns TO =1ns
.measure tran avgvall0bl263 AVG v(l0bl263) FROM = 0ns TO =1ns
.measure tran avgvall0bl264 AVG v(l0bl264) FROM = 0ns TO =1ns
.measure tran avgvall0bl265 AVG v(l0bl265) FROM = 0ns TO =1ns
.measure tran avgvall0bl266 AVG v(l0bl266) FROM = 0ns TO =1ns
.measure tran avgvall0bl267 AVG v(l0bl267) FROM = 0ns TO =1ns
.measure tran avgvall0bl268 AVG v(l0bl268) FROM = 0ns TO =1ns
.measure tran avgvall0bl269 AVG v(l0bl269) FROM = 0ns TO =1ns
.measure tran avgvall0bl270 AVG v(l0bl270) FROM = 0ns TO =1ns
.measure tran avgvall0bl271 AVG v(l0bl271) FROM = 0ns TO =1ns
.measure tran avgvall0bl272 AVG v(l0bl272) FROM = 0ns TO =1ns
.measure tran avgvall0bl273 AVG v(l0bl273) FROM = 0ns TO =1ns
.measure tran avgvall0bl274 AVG v(l0bl274) FROM = 0ns TO =1ns
.measure tran avgvall0bl275 AVG v(l0bl275) FROM = 0ns TO =1ns
.measure tran avgvall0bl276 AVG v(l0bl276) FROM = 0ns TO =1ns
.measure tran avgvall0bl277 AVG v(l0bl277) FROM = 0ns TO =1ns
.measure tran avgvall0bl278 AVG v(l0bl278) FROM = 0ns TO =1ns
.measure tran avgvall0bl279 AVG v(l0bl279) FROM = 0ns TO =1ns
.measure tran avgvall0bl280 AVG v(l0bl280) FROM = 0ns TO =1ns
.measure tran avgvall0bl281 AVG v(l0bl281) FROM = 0ns TO =1ns
.measure tran avgvall0bl282 AVG v(l0bl282) FROM = 0ns TO =1ns
.measure tran avgvall0bl283 AVG v(l0bl283) FROM = 0ns TO =1ns
.measure tran avgvall0bl284 AVG v(l0bl284) FROM = 0ns TO =1ns
.measure tran avgvall0bl285 AVG v(l0bl285) FROM = 0ns TO =1ns
.measure tran avgvall0bl286 AVG v(l0bl286) FROM = 0ns TO =1ns
.measure tran avgvall0bl287 AVG v(l0bl287) FROM = 0ns TO =1ns
.measure tran avgvall0bl288 AVG v(l0bl288) FROM = 0ns TO =1ns
.measure tran avgvall0bl289 AVG v(l0bl289) FROM = 0ns TO =1ns
.measure tran avgvall0bl290 AVG v(l0bl290) FROM = 0ns TO =1ns
.measure tran avgvall0bl291 AVG v(l0bl291) FROM = 0ns TO =1ns
.measure tran avgvall0bl292 AVG v(l0bl292) FROM = 0ns TO =1ns
.measure tran avgvall0bl293 AVG v(l0bl293) FROM = 0ns TO =1ns
.measure tran avgvall0bl294 AVG v(l0bl294) FROM = 0ns TO =1ns
.measure tran avgvall0bl295 AVG v(l0bl295) FROM = 0ns TO =1ns
.measure tran avgvall0bl296 AVG v(l0bl296) FROM = 0ns TO =1ns
.measure tran avgvall0bl297 AVG v(l0bl297) FROM = 0ns TO =1ns
.measure tran avgvall0bl298 AVG v(l0bl298) FROM = 0ns TO =1ns
.measure tran avgvall0bl299 AVG v(l0bl299) FROM = 0ns TO =1ns
.measure tran avgvall0bl300 AVG v(l0bl300) FROM = 0ns TO =1ns
.measure tran avgvall0bl301 AVG v(l0bl301) FROM = 0ns TO =1ns
.measure tran avgvall0bl302 AVG v(l0bl302) FROM = 0ns TO =1ns
.measure tran avgvall0bl303 AVG v(l0bl303) FROM = 0ns TO =1ns
.measure tran avgvall0bl304 AVG v(l0bl304) FROM = 0ns TO =1ns
.measure tran avgvall0bl305 AVG v(l0bl305) FROM = 0ns TO =1ns
.measure tran avgvall0bl306 AVG v(l0bl306) FROM = 0ns TO =1ns
.measure tran avgvall0bl307 AVG v(l0bl307) FROM = 0ns TO =1ns
.measure tran avgvall0bl308 AVG v(l0bl308) FROM = 0ns TO =1ns
.measure tran avgvall0bl309 AVG v(l0bl309) FROM = 0ns TO =1ns
.measure tran avgvall0bl310 AVG v(l0bl310) FROM = 0ns TO =1ns
.measure tran avgvall0bl311 AVG v(l0bl311) FROM = 0ns TO =1ns
.measure tran avgvall0bl312 AVG v(l0bl312) FROM = 0ns TO =1ns
.measure tran avgvall0bl313 AVG v(l0bl313) FROM = 0ns TO =1ns
.measure tran avgvall0bl314 AVG v(l0bl314) FROM = 0ns TO =1ns
.measure tran avgvall0bl315 AVG v(l0bl315) FROM = 0ns TO =1ns
.measure tran avgvall0bl316 AVG v(l0bl316) FROM = 0ns TO =1ns
.measure tran avgvall0bl317 AVG v(l0bl317) FROM = 0ns TO =1ns
.measure tran avgvall0bl318 AVG v(l0bl318) FROM = 0ns TO =1ns
.measure tran avgvall0bl319 AVG v(l0bl319) FROM = 0ns TO =1ns
.measure tran avgvall0bl320 AVG v(l0bl320) FROM = 0ns TO =1ns
.measure tran avgvall0bl321 AVG v(l0bl321) FROM = 0ns TO =1ns
.measure tran avgvall0bl322 AVG v(l0bl322) FROM = 0ns TO =1ns
.measure tran avgvall0bl323 AVG v(l0bl323) FROM = 0ns TO =1ns
.measure tran avgvall0bl324 AVG v(l0bl324) FROM = 0ns TO =1ns
.measure tran avgvall0bl325 AVG v(l0bl325) FROM = 0ns TO =1ns
.measure tran avgvall0bl326 AVG v(l0bl326) FROM = 0ns TO =1ns
.measure tran avgvall0bl327 AVG v(l0bl327) FROM = 0ns TO =1ns
.measure tran avgvall0bl328 AVG v(l0bl328) FROM = 0ns TO =1ns
.measure tran avgvall0bl329 AVG v(l0bl329) FROM = 0ns TO =1ns
.measure tran avgvall0bl330 AVG v(l0bl330) FROM = 0ns TO =1ns
.measure tran avgvall0bl331 AVG v(l0bl331) FROM = 0ns TO =1ns
.measure tran avgvall0bl332 AVG v(l0bl332) FROM = 0ns TO =1ns
.measure tran avgvall0bl333 AVG v(l0bl333) FROM = 0ns TO =1ns
.measure tran avgvall0bl334 AVG v(l0bl334) FROM = 0ns TO =1ns
.measure tran avgvall0bl335 AVG v(l0bl335) FROM = 0ns TO =1ns
.measure tran avgvall0bl336 AVG v(l0bl336) FROM = 0ns TO =1ns
.measure tran avgvall0bl337 AVG v(l0bl337) FROM = 0ns TO =1ns
.measure tran avgvall0bl338 AVG v(l0bl338) FROM = 0ns TO =1ns
.measure tran avgvall0bl339 AVG v(l0bl339) FROM = 0ns TO =1ns
.measure tran avgvall0bl340 AVG v(l0bl340) FROM = 0ns TO =1ns
.measure tran avgvall0bl341 AVG v(l0bl341) FROM = 0ns TO =1ns
.measure tran avgvall0bl342 AVG v(l0bl342) FROM = 0ns TO =1ns
.measure tran avgvall0bl343 AVG v(l0bl343) FROM = 0ns TO =1ns
.measure tran avgvall0bl344 AVG v(l0bl344) FROM = 0ns TO =1ns
.measure tran avgvall0bl345 AVG v(l0bl345) FROM = 0ns TO =1ns
.measure tran avgvall0bl346 AVG v(l0bl346) FROM = 0ns TO =1ns
.measure tran avgvall0bl347 AVG v(l0bl347) FROM = 0ns TO =1ns
.measure tran avgvall0bl348 AVG v(l0bl348) FROM = 0ns TO =1ns
.measure tran avgvall0bl349 AVG v(l0bl349) FROM = 0ns TO =1ns
.measure tran avgvall0bl350 AVG v(l0bl350) FROM = 0ns TO =1ns
.measure tran avgvall0bl351 AVG v(l0bl351) FROM = 0ns TO =1ns
.measure tran avgvall0bl352 AVG v(l0bl352) FROM = 0ns TO =1ns
.measure tran avgvall0bl353 AVG v(l0bl353) FROM = 0ns TO =1ns
.measure tran avgvall0bl354 AVG v(l0bl354) FROM = 0ns TO =1ns
.measure tran avgvall0bl355 AVG v(l0bl355) FROM = 0ns TO =1ns
.measure tran avgvall0bl356 AVG v(l0bl356) FROM = 0ns TO =1ns
.measure tran avgvall0bl357 AVG v(l0bl357) FROM = 0ns TO =1ns
.measure tran avgvall0bl358 AVG v(l0bl358) FROM = 0ns TO =1ns
.measure tran avgvall0bl359 AVG v(l0bl359) FROM = 0ns TO =1ns
.measure tran avgvall0bl360 AVG v(l0bl360) FROM = 0ns TO =1ns
.measure tran avgvall0bl361 AVG v(l0bl361) FROM = 0ns TO =1ns
.measure tran avgvall0bl362 AVG v(l0bl362) FROM = 0ns TO =1ns
.measure tran avgvall0bl363 AVG v(l0bl363) FROM = 0ns TO =1ns
.measure tran avgvall0bl364 AVG v(l0bl364) FROM = 0ns TO =1ns
.measure tran avgvall0bl365 AVG v(l0bl365) FROM = 0ns TO =1ns
.measure tran avgvall0bl366 AVG v(l0bl366) FROM = 0ns TO =1ns
.measure tran avgvall0bl367 AVG v(l0bl367) FROM = 0ns TO =1ns
.measure tran avgvall0bl368 AVG v(l0bl368) FROM = 0ns TO =1ns
.measure tran avgvall0bl369 AVG v(l0bl369) FROM = 0ns TO =1ns
.measure tran avgvall0bl370 AVG v(l0bl370) FROM = 0ns TO =1ns
.measure tran avgvall0bl371 AVG v(l0bl371) FROM = 0ns TO =1ns
.measure tran avgvall0bl372 AVG v(l0bl372) FROM = 0ns TO =1ns
.measure tran avgvall0bl373 AVG v(l0bl373) FROM = 0ns TO =1ns
.measure tran avgvall0bl374 AVG v(l0bl374) FROM = 0ns TO =1ns
.measure tran avgvall0bl375 AVG v(l0bl375) FROM = 0ns TO =1ns
.measure tran avgvall0bl376 AVG v(l0bl376) FROM = 0ns TO =1ns
.measure tran avgvall0bl377 AVG v(l0bl377) FROM = 0ns TO =1ns
.measure tran avgvall0bl378 AVG v(l0bl378) FROM = 0ns TO =1ns
.measure tran avgvall0bl379 AVG v(l0bl379) FROM = 0ns TO =1ns
.measure tran avgvall0bl380 AVG v(l0bl380) FROM = 0ns TO =1ns
.measure tran avgvall0bl381 AVG v(l0bl381) FROM = 0ns TO =1ns
.measure tran avgvall0bl382 AVG v(l0bl382) FROM = 0ns TO =1ns
.measure tran avgvall0bl383 AVG v(l0bl383) FROM = 0ns TO =1ns
.measure tran avgvall0bl384 AVG v(l0bl384) FROM = 0ns TO =1ns
.measure tran avgvall0bl385 AVG v(l0bl385) FROM = 0ns TO =1ns
.measure tran avgvall0bl386 AVG v(l0bl386) FROM = 0ns TO =1ns
.measure tran avgvall0bl387 AVG v(l0bl387) FROM = 0ns TO =1ns
.measure tran avgvall0bl388 AVG v(l0bl388) FROM = 0ns TO =1ns
.measure tran avgvall0bl389 AVG v(l0bl389) FROM = 0ns TO =1ns
.measure tran avgvall0bl390 AVG v(l0bl390) FROM = 0ns TO =1ns
.measure tran avgvall0bl391 AVG v(l0bl391) FROM = 0ns TO =1ns
.measure tran avgvall0bl392 AVG v(l0bl392) FROM = 0ns TO =1ns
.measure tran avgvall0bl393 AVG v(l0bl393) FROM = 0ns TO =1ns
.measure tran avgvall0bl394 AVG v(l0bl394) FROM = 0ns TO =1ns
.measure tran avgvall0bl395 AVG v(l0bl395) FROM = 0ns TO =1ns
.measure tran avgvall0bl396 AVG v(l0bl396) FROM = 0ns TO =1ns
.measure tran avgvall0bl397 AVG v(l0bl397) FROM = 0ns TO =1ns
.measure tran avgvall0bl398 AVG v(l0bl398) FROM = 0ns TO =1ns
.measure tran avgvall0bl399 AVG v(l0bl399) FROM = 0ns TO =1ns
.measure tran avgvall0bl400 AVG v(l0bl400) FROM = 0ns TO =1ns
.measure tran avgvall0bl401 AVG v(l0bl401) FROM = 0ns TO =1ns
.measure tran avgvall0bl402 AVG v(l0bl402) FROM = 0ns TO =1ns
.measure tran avgvall0bl403 AVG v(l0bl403) FROM = 0ns TO =1ns
.measure tran avgvall0bl404 AVG v(l0bl404) FROM = 0ns TO =1ns
.measure tran avgvall0bl405 AVG v(l0bl405) FROM = 0ns TO =1ns
.measure tran avgvall0bl406 AVG v(l0bl406) FROM = 0ns TO =1ns
.measure tran avgvall0bl407 AVG v(l0bl407) FROM = 0ns TO =1ns
.measure tran avgvall0bl408 AVG v(l0bl408) FROM = 0ns TO =1ns
.measure tran avgvall0bl409 AVG v(l0bl409) FROM = 0ns TO =1ns
.measure tran avgvall0bl410 AVG v(l0bl410) FROM = 0ns TO =1ns
.measure tran avgvall0bl411 AVG v(l0bl411) FROM = 0ns TO =1ns
.measure tran avgvall0bl412 AVG v(l0bl412) FROM = 0ns TO =1ns
.measure tran avgvall0bl413 AVG v(l0bl413) FROM = 0ns TO =1ns
.measure tran avgvall0bl414 AVG v(l0bl414) FROM = 0ns TO =1ns
.measure tran avgvall0bl415 AVG v(l0bl415) FROM = 0ns TO =1ns
.measure tran avgvall0bl416 AVG v(l0bl416) FROM = 0ns TO =1ns
.measure tran avgvall0bl417 AVG v(l0bl417) FROM = 0ns TO =1ns
.measure tran avgvall0bl418 AVG v(l0bl418) FROM = 0ns TO =1ns
.measure tran avgvall0bl419 AVG v(l0bl419) FROM = 0ns TO =1ns
.measure tran avgvall0bl420 AVG v(l0bl420) FROM = 0ns TO =1ns
.measure tran avgvall0bl421 AVG v(l0bl421) FROM = 0ns TO =1ns
.measure tran avgvall0bl422 AVG v(l0bl422) FROM = 0ns TO =1ns
.measure tran avgvall0bl423 AVG v(l0bl423) FROM = 0ns TO =1ns
.measure tran avgvall0bl424 AVG v(l0bl424) FROM = 0ns TO =1ns
.measure tran avgvall0bl425 AVG v(l0bl425) FROM = 0ns TO =1ns
.measure tran avgvall0bl426 AVG v(l0bl426) FROM = 0ns TO =1ns
.measure tran avgvall0bl427 AVG v(l0bl427) FROM = 0ns TO =1ns
.measure tran avgvall0bl428 AVG v(l0bl428) FROM = 0ns TO =1ns
.measure tran avgvall0bl429 AVG v(l0bl429) FROM = 0ns TO =1ns
.measure tran avgvall0bl430 AVG v(l0bl430) FROM = 0ns TO =1ns
.measure tran avgvall0bl431 AVG v(l0bl431) FROM = 0ns TO =1ns
.measure tran avgvall0bl432 AVG v(l0bl432) FROM = 0ns TO =1ns
.measure tran avgvall0bl433 AVG v(l0bl433) FROM = 0ns TO =1ns
.measure tran avgvall0bl434 AVG v(l0bl434) FROM = 0ns TO =1ns
.measure tran avgvall0bl435 AVG v(l0bl435) FROM = 0ns TO =1ns
.measure tran avgvall0bl436 AVG v(l0bl436) FROM = 0ns TO =1ns
.measure tran avgvall0bl437 AVG v(l0bl437) FROM = 0ns TO =1ns
.measure tran avgvall0bl438 AVG v(l0bl438) FROM = 0ns TO =1ns
.measure tran avgvall0bl439 AVG v(l0bl439) FROM = 0ns TO =1ns
.measure tran avgvall0bl440 AVG v(l0bl440) FROM = 0ns TO =1ns
.measure tran avgvall0bl441 AVG v(l0bl441) FROM = 0ns TO =1ns
.measure tran avgvall0bl442 AVG v(l0bl442) FROM = 0ns TO =1ns
.measure tran avgvall0bl443 AVG v(l0bl443) FROM = 0ns TO =1ns
.measure tran avgvall0bl444 AVG v(l0bl444) FROM = 0ns TO =1ns
.measure tran avgvall0bl445 AVG v(l0bl445) FROM = 0ns TO =1ns
.measure tran avgvall0bl446 AVG v(l0bl446) FROM = 0ns TO =1ns
.measure tran avgvall0bl447 AVG v(l0bl447) FROM = 0ns TO =1ns
.measure tran avgvall0bl448 AVG v(l0bl448) FROM = 0ns TO =1ns
.measure tran avgvall0bl449 AVG v(l0bl449) FROM = 0ns TO =1ns
.measure tran avgvall0bl450 AVG v(l0bl450) FROM = 0ns TO =1ns
.measure tran avgvall0bl451 AVG v(l0bl451) FROM = 0ns TO =1ns
.measure tran avgvall0bl452 AVG v(l0bl452) FROM = 0ns TO =1ns
.measure tran avgvall0bl453 AVG v(l0bl453) FROM = 0ns TO =1ns
.measure tran avgvall0bl454 AVG v(l0bl454) FROM = 0ns TO =1ns
.measure tran avgvall0bl455 AVG v(l0bl455) FROM = 0ns TO =1ns
.measure tran avgvall0bl456 AVG v(l0bl456) FROM = 0ns TO =1ns
.measure tran avgvall0bl457 AVG v(l0bl457) FROM = 0ns TO =1ns
.measure tran avgvall0bl458 AVG v(l0bl458) FROM = 0ns TO =1ns
.measure tran avgvall0bl459 AVG v(l0bl459) FROM = 0ns TO =1ns
.measure tran avgvall0bl460 AVG v(l0bl460) FROM = 0ns TO =1ns
.measure tran avgvall0bl461 AVG v(l0bl461) FROM = 0ns TO =1ns
.measure tran avgvall0bl462 AVG v(l0bl462) FROM = 0ns TO =1ns
.measure tran avgvall0bl463 AVG v(l0bl463) FROM = 0ns TO =1ns
.measure tran avgvall0bl464 AVG v(l0bl464) FROM = 0ns TO =1ns
.measure tran avgvall0bl465 AVG v(l0bl465) FROM = 0ns TO =1ns
.measure tran avgvall0bl466 AVG v(l0bl466) FROM = 0ns TO =1ns
.measure tran avgvall0bl467 AVG v(l0bl467) FROM = 0ns TO =1ns
.measure tran avgvall0bl468 AVG v(l0bl468) FROM = 0ns TO =1ns
.measure tran avgvall0bl469 AVG v(l0bl469) FROM = 0ns TO =1ns
.measure tran avgvall0bl470 AVG v(l0bl470) FROM = 0ns TO =1ns
.measure tran avgvall0bl471 AVG v(l0bl471) FROM = 0ns TO =1ns
.measure tran avgvall0bl472 AVG v(l0bl472) FROM = 0ns TO =1ns
.measure tran avgvall0bl473 AVG v(l0bl473) FROM = 0ns TO =1ns
.measure tran avgvall0bl474 AVG v(l0bl474) FROM = 0ns TO =1ns
.measure tran avgvall0bl475 AVG v(l0bl475) FROM = 0ns TO =1ns
.measure tran avgvall0bl476 AVG v(l0bl476) FROM = 0ns TO =1ns
.measure tran avgvall0bl477 AVG v(l0bl477) FROM = 0ns TO =1ns
.measure tran avgvall0bl478 AVG v(l0bl478) FROM = 0ns TO =1ns
.measure tran avgvall0bl479 AVG v(l0bl479) FROM = 0ns TO =1ns
.measure tran avgvall0bl480 AVG v(l0bl480) FROM = 0ns TO =1ns
.measure tran avgvall0bl481 AVG v(l0bl481) FROM = 0ns TO =1ns
.measure tran avgvall0bl482 AVG v(l0bl482) FROM = 0ns TO =1ns
.measure tran avgvall0bl483 AVG v(l0bl483) FROM = 0ns TO =1ns
.measure tran avgvall0bl484 AVG v(l0bl484) FROM = 0ns TO =1ns
.measure tran avgvall0bl485 AVG v(l0bl485) FROM = 0ns TO =1ns
.measure tran avgvall0bl486 AVG v(l0bl486) FROM = 0ns TO =1ns
.measure tran avgvall0bl487 AVG v(l0bl487) FROM = 0ns TO =1ns
.measure tran avgvall0bl488 AVG v(l0bl488) FROM = 0ns TO =1ns
.measure tran avgvall0bl489 AVG v(l0bl489) FROM = 0ns TO =1ns
.measure tran avgvall0bl490 AVG v(l0bl490) FROM = 0ns TO =1ns
.measure tran avgvall0bl491 AVG v(l0bl491) FROM = 0ns TO =1ns
.measure tran avgvall0bl492 AVG v(l0bl492) FROM = 0ns TO =1ns
.measure tran avgvall0bl493 AVG v(l0bl493) FROM = 0ns TO =1ns
.measure tran avgvall0bl494 AVG v(l0bl494) FROM = 0ns TO =1ns
.measure tran avgvall0bl495 AVG v(l0bl495) FROM = 0ns TO =1ns
.measure tran avgvall0bl496 AVG v(l0bl496) FROM = 0ns TO =1ns
.measure tran avgvall0bl497 AVG v(l0bl497) FROM = 0ns TO =1ns
.measure tran avgvall0bl498 AVG v(l0bl498) FROM = 0ns TO =1ns
.measure tran avgvall0bl499 AVG v(l0bl499) FROM = 0ns TO =1ns
.measure tran avgvall0bl500 AVG v(l0bl500) FROM = 0ns TO =1ns
.measure tran avgvall0bl501 AVG v(l0bl501) FROM = 0ns TO =1ns
.measure tran avgvall0bl502 AVG v(l0bl502) FROM = 0ns TO =1ns
.measure tran avgvall0bl503 AVG v(l0bl503) FROM = 0ns TO =1ns
.measure tran avgvall0bl504 AVG v(l0bl504) FROM = 0ns TO =1ns
.measure tran avgvall0bl505 AVG v(l0bl505) FROM = 0ns TO =1ns
.measure tran avgvall0bl506 AVG v(l0bl506) FROM = 0ns TO =1ns
.measure tran avgvall0bl507 AVG v(l0bl507) FROM = 0ns TO =1ns
.measure tran avgvall0bl508 AVG v(l0bl508) FROM = 0ns TO =1ns
.measure tran avgvall0bl509 AVG v(l0bl509) FROM = 0ns TO =1ns
.measure tran avgvall0bl510 AVG v(l0bl510) FROM = 0ns TO =1ns
.measure tran avgvall0bl511 AVG v(l0bl511) FROM = 0ns TO =1ns

.measure tran avgvall1bl0 AVG v(l1bl0) FROM = 199ns TO =200ns
.measure tran avgvall1bl1 AVG v(l1bl1) FROM = 199ns TO =200ns
.measure tran avgvall1bl2 AVG v(l1bl2) FROM = 199ns TO =200ns
.measure tran avgvall1bl3 AVG v(l1bl3) FROM = 199ns TO =200ns
.measure tran avgvall1bl4 AVG v(l1bl4) FROM = 199ns TO =200ns
.measure tran avgvall1bl5 AVG v(l1bl5) FROM = 199ns TO =200ns
.measure tran avgvall1bl6 AVG v(l1bl6) FROM = 199ns TO =200ns
.measure tran avgvall1bl7 AVG v(l1bl7) FROM = 199ns TO =200ns
.measure tran avgvall1bl8 AVG v(l1bl8) FROM = 199ns TO =200ns
.measure tran avgvall1bl9 AVG v(l1bl9) FROM = 199ns TO =200ns
.measure tran avgvall1bl10 AVG v(l1bl10) FROM = 199ns TO =200ns
.measure tran avgvall1bl11 AVG v(l1bl11) FROM = 199ns TO =200ns
.measure tran avgvall1bl12 AVG v(l1bl12) FROM = 199ns TO =200ns
.measure tran avgvall1bl13 AVG v(l1bl13) FROM = 199ns TO =200ns
.measure tran avgvall1bl14 AVG v(l1bl14) FROM = 199ns TO =200ns
.measure tran avgvall1bl15 AVG v(l1bl15) FROM = 199ns TO =200ns
.measure tran avgvall1bl16 AVG v(l1bl16) FROM = 199ns TO =200ns
.measure tran avgvall1bl17 AVG v(l1bl17) FROM = 199ns TO =200ns
.measure tran avgvall1bl18 AVG v(l1bl18) FROM = 199ns TO =200ns
.measure tran avgvall1bl19 AVG v(l1bl19) FROM = 199ns TO =200ns
.measure tran avgvall1bl20 AVG v(l1bl20) FROM = 199ns TO =200ns
.measure tran avgvall1bl21 AVG v(l1bl21) FROM = 199ns TO =200ns
.measure tran avgvall1bl22 AVG v(l1bl22) FROM = 199ns TO =200ns
.measure tran avgvall1bl23 AVG v(l1bl23) FROM = 199ns TO =200ns
.measure tran avgvall1bl24 AVG v(l1bl24) FROM = 199ns TO =200ns
.measure tran avgvall1bl25 AVG v(l1bl25) FROM = 199ns TO =200ns
.measure tran avgvall1bl26 AVG v(l1bl26) FROM = 199ns TO =200ns
.measure tran avgvall1bl27 AVG v(l1bl27) FROM = 199ns TO =200ns
.measure tran avgvall1bl28 AVG v(l1bl28) FROM = 199ns TO =200ns
.measure tran avgvall1bl29 AVG v(l1bl29) FROM = 199ns TO =200ns
.measure tran avgvall1bl30 AVG v(l1bl30) FROM = 199ns TO =200ns
.measure tran avgvall1bl31 AVG v(l1bl31) FROM = 199ns TO =200ns
.measure tran avgvall1bl32 AVG v(l1bl32) FROM = 199ns TO =200ns
.measure tran avgvall1bl33 AVG v(l1bl33) FROM = 199ns TO =200ns
.measure tran avgvall1bl34 AVG v(l1bl34) FROM = 199ns TO =200ns
.measure tran avgvall1bl35 AVG v(l1bl35) FROM = 199ns TO =200ns
.measure tran avgvall1bl36 AVG v(l1bl36) FROM = 199ns TO =200ns
.measure tran avgvall1bl37 AVG v(l1bl37) FROM = 199ns TO =200ns
.measure tran avgvall1bl38 AVG v(l1bl38) FROM = 199ns TO =200ns
.measure tran avgvall1bl39 AVG v(l1bl39) FROM = 199ns TO =200ns
.measure tran avgvall1bl40 AVG v(l1bl40) FROM = 199ns TO =200ns
.measure tran avgvall1bl41 AVG v(l1bl41) FROM = 199ns TO =200ns
.measure tran avgvall1bl42 AVG v(l1bl42) FROM = 199ns TO =200ns
.measure tran avgvall1bl43 AVG v(l1bl43) FROM = 199ns TO =200ns
.measure tran avgvall1bl44 AVG v(l1bl44) FROM = 199ns TO =200ns
.measure tran avgvall1bl45 AVG v(l1bl45) FROM = 199ns TO =200ns
.measure tran avgvall1bl46 AVG v(l1bl46) FROM = 199ns TO =200ns
.measure tran avgvall1bl47 AVG v(l1bl47) FROM = 199ns TO =200ns
.measure tran avgvall1bl48 AVG v(l1bl48) FROM = 199ns TO =200ns
.measure tran avgvall1bl49 AVG v(l1bl49) FROM = 199ns TO =200ns
.measure tran avgvall1bl50 AVG v(l1bl50) FROM = 199ns TO =200ns
.measure tran avgvall1bl51 AVG v(l1bl51) FROM = 199ns TO =200ns
.measure tran avgvall1bl52 AVG v(l1bl52) FROM = 199ns TO =200ns
.measure tran avgvall1bl53 AVG v(l1bl53) FROM = 199ns TO =200ns
.measure tran avgvall1bl54 AVG v(l1bl54) FROM = 199ns TO =200ns
.measure tran avgvall1bl55 AVG v(l1bl55) FROM = 199ns TO =200ns
.measure tran avgvall1bl56 AVG v(l1bl56) FROM = 199ns TO =200ns
.measure tran avgvall1bl57 AVG v(l1bl57) FROM = 199ns TO =200ns
.measure tran avgvall1bl58 AVG v(l1bl58) FROM = 199ns TO =200ns
.measure tran avgvall1bl59 AVG v(l1bl59) FROM = 199ns TO =200ns
.measure tran avgvall1bl60 AVG v(l1bl60) FROM = 199ns TO =200ns
.measure tran avgvall1bl61 AVG v(l1bl61) FROM = 199ns TO =200ns
.measure tran avgvall1bl62 AVG v(l1bl62) FROM = 199ns TO =200ns
.measure tran avgvall1bl63 AVG v(l1bl63) FROM = 199ns TO =200ns
.measure tran avgvall1bl64 AVG v(l1bl64) FROM = 199ns TO =200ns
.measure tran avgvall1bl65 AVG v(l1bl65) FROM = 199ns TO =200ns
.measure tran avgvall1bl66 AVG v(l1bl66) FROM = 199ns TO =200ns
.measure tran avgvall1bl67 AVG v(l1bl67) FROM = 199ns TO =200ns
.measure tran avgvall1bl68 AVG v(l1bl68) FROM = 199ns TO =200ns
.measure tran avgvall1bl69 AVG v(l1bl69) FROM = 199ns TO =200ns
.measure tran avgvall1bl70 AVG v(l1bl70) FROM = 199ns TO =200ns
.measure tran avgvall1bl71 AVG v(l1bl71) FROM = 199ns TO =200ns
.measure tran avgvall1bl72 AVG v(l1bl72) FROM = 199ns TO =200ns
.measure tran avgvall1bl73 AVG v(l1bl73) FROM = 199ns TO =200ns
.measure tran avgvall1bl74 AVG v(l1bl74) FROM = 199ns TO =200ns
.measure tran avgvall1bl75 AVG v(l1bl75) FROM = 199ns TO =200ns
.measure tran avgvall1bl76 AVG v(l1bl76) FROM = 199ns TO =200ns
.measure tran avgvall1bl77 AVG v(l1bl77) FROM = 199ns TO =200ns
.measure tran avgvall1bl78 AVG v(l1bl78) FROM = 199ns TO =200ns
.measure tran avgvall1bl79 AVG v(l1bl79) FROM = 199ns TO =200ns
.measure tran avgvall1bl80 AVG v(l1bl80) FROM = 199ns TO =200ns
.measure tran avgvall1bl81 AVG v(l1bl81) FROM = 199ns TO =200ns
.measure tran avgvall1bl82 AVG v(l1bl82) FROM = 199ns TO =200ns
.measure tran avgvall1bl83 AVG v(l1bl83) FROM = 199ns TO =200ns
.measure tran avgvall1bl84 AVG v(l1bl84) FROM = 199ns TO =200ns
.measure tran avgvall1bl85 AVG v(l1bl85) FROM = 199ns TO =200ns
.measure tran avgvall1bl86 AVG v(l1bl86) FROM = 199ns TO =200ns
.measure tran avgvall1bl87 AVG v(l1bl87) FROM = 199ns TO =200ns
.measure tran avgvall1bl88 AVG v(l1bl88) FROM = 199ns TO =200ns
.measure tran avgvall1bl89 AVG v(l1bl89) FROM = 199ns TO =200ns
.measure tran avgvall1bl90 AVG v(l1bl90) FROM = 199ns TO =200ns
.measure tran avgvall1bl91 AVG v(l1bl91) FROM = 199ns TO =200ns
.measure tran avgvall1bl92 AVG v(l1bl92) FROM = 199ns TO =200ns
.measure tran avgvall1bl93 AVG v(l1bl93) FROM = 199ns TO =200ns
.measure tran avgvall1bl94 AVG v(l1bl94) FROM = 199ns TO =200ns
.measure tran avgvall1bl95 AVG v(l1bl95) FROM = 199ns TO =200ns
.measure tran avgvall1bl96 AVG v(l1bl96) FROM = 199ns TO =200ns
.measure tran avgvall1bl97 AVG v(l1bl97) FROM = 199ns TO =200ns
.measure tran avgvall1bl98 AVG v(l1bl98) FROM = 199ns TO =200ns
.measure tran avgvall1bl99 AVG v(l1bl99) FROM = 199ns TO =200ns
.measure tran avgvall1bl100 AVG v(l1bl100) FROM = 199ns TO =200ns
.measure tran avgvall1bl101 AVG v(l1bl101) FROM = 199ns TO =200ns
.measure tran avgvall1bl102 AVG v(l1bl102) FROM = 199ns TO =200ns
.measure tran avgvall1bl103 AVG v(l1bl103) FROM = 199ns TO =200ns
.measure tran avgvall1bl104 AVG v(l1bl104) FROM = 199ns TO =200ns
.measure tran avgvall1bl105 AVG v(l1bl105) FROM = 199ns TO =200ns
.measure tran avgvall1bl106 AVG v(l1bl106) FROM = 199ns TO =200ns
.measure tran avgvall1bl107 AVG v(l1bl107) FROM = 199ns TO =200ns
.measure tran avgvall1bl108 AVG v(l1bl108) FROM = 199ns TO =200ns
.measure tran avgvall1bl109 AVG v(l1bl109) FROM = 199ns TO =200ns
.measure tran avgvall1bl110 AVG v(l1bl110) FROM = 199ns TO =200ns
.measure tran avgvall1bl111 AVG v(l1bl111) FROM = 199ns TO =200ns
.measure tran avgvall1bl112 AVG v(l1bl112) FROM = 199ns TO =200ns
.measure tran avgvall1bl113 AVG v(l1bl113) FROM = 199ns TO =200ns
.measure tran avgvall1bl114 AVG v(l1bl114) FROM = 199ns TO =200ns
.measure tran avgvall1bl115 AVG v(l1bl115) FROM = 199ns TO =200ns
.measure tran avgvall1bl116 AVG v(l1bl116) FROM = 199ns TO =200ns
.measure tran avgvall1bl117 AVG v(l1bl117) FROM = 199ns TO =200ns
.measure tran avgvall1bl118 AVG v(l1bl118) FROM = 199ns TO =200ns
.measure tran avgvall1bl119 AVG v(l1bl119) FROM = 199ns TO =200ns
.measure tran avgvall1bl120 AVG v(l1bl120) FROM = 199ns TO =200ns
.measure tran avgvall1bl121 AVG v(l1bl121) FROM = 199ns TO =200ns
.measure tran avgvall1bl122 AVG v(l1bl122) FROM = 199ns TO =200ns
.measure tran avgvall1bl123 AVG v(l1bl123) FROM = 199ns TO =200ns
.measure tran avgvall1bl124 AVG v(l1bl124) FROM = 199ns TO =200ns
.measure tran avgvall1bl125 AVG v(l1bl125) FROM = 199ns TO =200ns
.measure tran avgvall1bl126 AVG v(l1bl126) FROM = 199ns TO =200ns
.measure tran avgvall1bl127 AVG v(l1bl127) FROM = 199ns TO =200ns
.measure tran avgvall1bl128 AVG v(l1bl128) FROM = 199ns TO =200ns
.measure tran avgvall1bl129 AVG v(l1bl129) FROM = 199ns TO =200ns
.measure tran avgvall1bl130 AVG v(l1bl130) FROM = 199ns TO =200ns
.measure tran avgvall1bl131 AVG v(l1bl131) FROM = 199ns TO =200ns
.measure tran avgvall1bl132 AVG v(l1bl132) FROM = 199ns TO =200ns
.measure tran avgvall1bl133 AVG v(l1bl133) FROM = 199ns TO =200ns
.measure tran avgvall1bl134 AVG v(l1bl134) FROM = 199ns TO =200ns
.measure tran avgvall1bl135 AVG v(l1bl135) FROM = 199ns TO =200ns
.measure tran avgvall1bl136 AVG v(l1bl136) FROM = 199ns TO =200ns
.measure tran avgvall1bl137 AVG v(l1bl137) FROM = 199ns TO =200ns
.measure tran avgvall1bl138 AVG v(l1bl138) FROM = 199ns TO =200ns
.measure tran avgvall1bl139 AVG v(l1bl139) FROM = 199ns TO =200ns
.measure tran avgvall1bl140 AVG v(l1bl140) FROM = 199ns TO =200ns
.measure tran avgvall1bl141 AVG v(l1bl141) FROM = 199ns TO =200ns
.measure tran avgvall1bl142 AVG v(l1bl142) FROM = 199ns TO =200ns
.measure tran avgvall1bl143 AVG v(l1bl143) FROM = 199ns TO =200ns
.measure tran avgvall1bl144 AVG v(l1bl144) FROM = 199ns TO =200ns
.measure tran avgvall1bl145 AVG v(l1bl145) FROM = 199ns TO =200ns
.measure tran avgvall1bl146 AVG v(l1bl146) FROM = 199ns TO =200ns
.measure tran avgvall1bl147 AVG v(l1bl147) FROM = 199ns TO =200ns
.measure tran avgvall1bl148 AVG v(l1bl148) FROM = 199ns TO =200ns
.measure tran avgvall1bl149 AVG v(l1bl149) FROM = 199ns TO =200ns
.measure tran avgvall1bl150 AVG v(l1bl150) FROM = 199ns TO =200ns
.measure tran avgvall1bl151 AVG v(l1bl151) FROM = 199ns TO =200ns
.measure tran avgvall1bl152 AVG v(l1bl152) FROM = 199ns TO =200ns
.measure tran avgvall1bl153 AVG v(l1bl153) FROM = 199ns TO =200ns
.measure tran avgvall1bl154 AVG v(l1bl154) FROM = 199ns TO =200ns
.measure tran avgvall1bl155 AVG v(l1bl155) FROM = 199ns TO =200ns
.measure tran avgvall1bl156 AVG v(l1bl156) FROM = 199ns TO =200ns
.measure tran avgvall1bl157 AVG v(l1bl157) FROM = 199ns TO =200ns
.measure tran avgvall1bl158 AVG v(l1bl158) FROM = 199ns TO =200ns
.measure tran avgvall1bl159 AVG v(l1bl159) FROM = 199ns TO =200ns
.measure tran avgvall1bl160 AVG v(l1bl160) FROM = 199ns TO =200ns
.measure tran avgvall1bl161 AVG v(l1bl161) FROM = 199ns TO =200ns
.measure tran avgvall1bl162 AVG v(l1bl162) FROM = 199ns TO =200ns
.measure tran avgvall1bl163 AVG v(l1bl163) FROM = 199ns TO =200ns
.measure tran avgvall1bl164 AVG v(l1bl164) FROM = 199ns TO =200ns
.measure tran avgvall1bl165 AVG v(l1bl165) FROM = 199ns TO =200ns
.measure tran avgvall1bl166 AVG v(l1bl166) FROM = 199ns TO =200ns
.measure tran avgvall1bl167 AVG v(l1bl167) FROM = 199ns TO =200ns
.measure tran avgvall1bl168 AVG v(l1bl168) FROM = 199ns TO =200ns
.measure tran avgvall1bl169 AVG v(l1bl169) FROM = 199ns TO =200ns
.measure tran avgvall1bl170 AVG v(l1bl170) FROM = 199ns TO =200ns
.measure tran avgvall1bl171 AVG v(l1bl171) FROM = 199ns TO =200ns
.measure tran avgvall1bl172 AVG v(l1bl172) FROM = 199ns TO =200ns
.measure tran avgvall1bl173 AVG v(l1bl173) FROM = 199ns TO =200ns
.measure tran avgvall1bl174 AVG v(l1bl174) FROM = 199ns TO =200ns
.measure tran avgvall1bl175 AVG v(l1bl175) FROM = 199ns TO =200ns
.measure tran avgvall1bl176 AVG v(l1bl176) FROM = 199ns TO =200ns
.measure tran avgvall1bl177 AVG v(l1bl177) FROM = 199ns TO =200ns
.measure tran avgvall1bl178 AVG v(l1bl178) FROM = 199ns TO =200ns
.measure tran avgvall1bl179 AVG v(l1bl179) FROM = 199ns TO =200ns
.measure tran avgvall1bl180 AVG v(l1bl180) FROM = 199ns TO =200ns
.measure tran avgvall1bl181 AVG v(l1bl181) FROM = 199ns TO =200ns
.measure tran avgvall1bl182 AVG v(l1bl182) FROM = 199ns TO =200ns
.measure tran avgvall1bl183 AVG v(l1bl183) FROM = 199ns TO =200ns
.measure tran avgvall1bl184 AVG v(l1bl184) FROM = 199ns TO =200ns
.measure tran avgvall1bl185 AVG v(l1bl185) FROM = 199ns TO =200ns
.measure tran avgvall1bl186 AVG v(l1bl186) FROM = 199ns TO =200ns
.measure tran avgvall1bl187 AVG v(l1bl187) FROM = 199ns TO =200ns
.measure tran avgvall1bl188 AVG v(l1bl188) FROM = 199ns TO =200ns
.measure tran avgvall1bl189 AVG v(l1bl189) FROM = 199ns TO =200ns
.measure tran avgvall1bl190 AVG v(l1bl190) FROM = 199ns TO =200ns
.measure tran avgvall1bl191 AVG v(l1bl191) FROM = 199ns TO =200ns
.measure tran avgvall1bl192 AVG v(l1bl192) FROM = 199ns TO =200ns
.measure tran avgvall1bl193 AVG v(l1bl193) FROM = 199ns TO =200ns
.measure tran avgvall1bl194 AVG v(l1bl194) FROM = 199ns TO =200ns
.measure tran avgvall1bl195 AVG v(l1bl195) FROM = 199ns TO =200ns
.measure tran avgvall1bl196 AVG v(l1bl196) FROM = 199ns TO =200ns
.measure tran avgvall1bl197 AVG v(l1bl197) FROM = 199ns TO =200ns
.measure tran avgvall1bl198 AVG v(l1bl198) FROM = 199ns TO =200ns
.measure tran avgvall1bl199 AVG v(l1bl199) FROM = 199ns TO =200ns
.measure tran avgvall1bl200 AVG v(l1bl200) FROM = 199ns TO =200ns
.measure tran avgvall1bl201 AVG v(l1bl201) FROM = 199ns TO =200ns
.measure tran avgvall1bl202 AVG v(l1bl202) FROM = 199ns TO =200ns
.measure tran avgvall1bl203 AVG v(l1bl203) FROM = 199ns TO =200ns
.measure tran avgvall1bl204 AVG v(l1bl204) FROM = 199ns TO =200ns
.measure tran avgvall1bl205 AVG v(l1bl205) FROM = 199ns TO =200ns
.measure tran avgvall1bl206 AVG v(l1bl206) FROM = 199ns TO =200ns
.measure tran avgvall1bl207 AVG v(l1bl207) FROM = 199ns TO =200ns
.measure tran avgvall1bl208 AVG v(l1bl208) FROM = 199ns TO =200ns
.measure tran avgvall1bl209 AVG v(l1bl209) FROM = 199ns TO =200ns
.measure tran avgvall1bl210 AVG v(l1bl210) FROM = 199ns TO =200ns
.measure tran avgvall1bl211 AVG v(l1bl211) FROM = 199ns TO =200ns
.measure tran avgvall1bl212 AVG v(l1bl212) FROM = 199ns TO =200ns
.measure tran avgvall1bl213 AVG v(l1bl213) FROM = 199ns TO =200ns
.measure tran avgvall1bl214 AVG v(l1bl214) FROM = 199ns TO =200ns
.measure tran avgvall1bl215 AVG v(l1bl215) FROM = 199ns TO =200ns
.measure tran avgvall1bl216 AVG v(l1bl216) FROM = 199ns TO =200ns
.measure tran avgvall1bl217 AVG v(l1bl217) FROM = 199ns TO =200ns
.measure tran avgvall1bl218 AVG v(l1bl218) FROM = 199ns TO =200ns
.measure tran avgvall1bl219 AVG v(l1bl219) FROM = 199ns TO =200ns
.measure tran avgvall1bl220 AVG v(l1bl220) FROM = 199ns TO =200ns
.measure tran avgvall1bl221 AVG v(l1bl221) FROM = 199ns TO =200ns
.measure tran avgvall1bl222 AVG v(l1bl222) FROM = 199ns TO =200ns
.measure tran avgvall1bl223 AVG v(l1bl223) FROM = 199ns TO =200ns
.measure tran avgvall1bl224 AVG v(l1bl224) FROM = 199ns TO =200ns
.measure tran avgvall1bl225 AVG v(l1bl225) FROM = 199ns TO =200ns
.measure tran avgvall1bl226 AVG v(l1bl226) FROM = 199ns TO =200ns
.measure tran avgvall1bl227 AVG v(l1bl227) FROM = 199ns TO =200ns
.measure tran avgvall1bl228 AVG v(l1bl228) FROM = 199ns TO =200ns
.measure tran avgvall1bl229 AVG v(l1bl229) FROM = 199ns TO =200ns
.measure tran avgvall1bl230 AVG v(l1bl230) FROM = 199ns TO =200ns
.measure tran avgvall1bl231 AVG v(l1bl231) FROM = 199ns TO =200ns
.measure tran avgvall1bl232 AVG v(l1bl232) FROM = 199ns TO =200ns
.measure tran avgvall1bl233 AVG v(l1bl233) FROM = 199ns TO =200ns
.measure tran avgvall1bl234 AVG v(l1bl234) FROM = 199ns TO =200ns
.measure tran avgvall1bl235 AVG v(l1bl235) FROM = 199ns TO =200ns
.measure tran avgvall1bl236 AVG v(l1bl236) FROM = 199ns TO =200ns
.measure tran avgvall1bl237 AVG v(l1bl237) FROM = 199ns TO =200ns
.measure tran avgvall1bl238 AVG v(l1bl238) FROM = 199ns TO =200ns
.measure tran avgvall1bl239 AVG v(l1bl239) FROM = 199ns TO =200ns
.measure tran avgvall1bl240 AVG v(l1bl240) FROM = 199ns TO =200ns
.measure tran avgvall1bl241 AVG v(l1bl241) FROM = 199ns TO =200ns
.measure tran avgvall1bl242 AVG v(l1bl242) FROM = 199ns TO =200ns
.measure tran avgvall1bl243 AVG v(l1bl243) FROM = 199ns TO =200ns
.measure tran avgvall1bl244 AVG v(l1bl244) FROM = 199ns TO =200ns
.measure tran avgvall1bl245 AVG v(l1bl245) FROM = 199ns TO =200ns
.measure tran avgvall1bl246 AVG v(l1bl246) FROM = 199ns TO =200ns
.measure tran avgvall1bl247 AVG v(l1bl247) FROM = 199ns TO =200ns
.measure tran avgvall1bl248 AVG v(l1bl248) FROM = 199ns TO =200ns
.measure tran avgvall1bl249 AVG v(l1bl249) FROM = 199ns TO =200ns
.measure tran avgvall1bl250 AVG v(l1bl250) FROM = 199ns TO =200ns
.measure tran avgvall1bl251 AVG v(l1bl251) FROM = 199ns TO =200ns
.measure tran avgvall1bl252 AVG v(l1bl252) FROM = 199ns TO =200ns
.measure tran avgvall1bl253 AVG v(l1bl253) FROM = 199ns TO =200ns
.measure tran avgvall1bl254 AVG v(l1bl254) FROM = 199ns TO =200ns
.measure tran avgvall1bl255 AVG v(l1bl255) FROM = 199ns TO =200ns
.measure tran avgvall1bl256 AVG v(l1bl256) FROM = 199ns TO =200ns
.measure tran avgvall1bl257 AVG v(l1bl257) FROM = 199ns TO =200ns
.measure tran avgvall1bl258 AVG v(l1bl258) FROM = 199ns TO =200ns
.measure tran avgvall1bl259 AVG v(l1bl259) FROM = 199ns TO =200ns
.measure tran avgvall1bl260 AVG v(l1bl260) FROM = 199ns TO =200ns
.measure tran avgvall1bl261 AVG v(l1bl261) FROM = 199ns TO =200ns
.measure tran avgvall1bl262 AVG v(l1bl262) FROM = 199ns TO =200ns
.measure tran avgvall1bl263 AVG v(l1bl263) FROM = 199ns TO =200ns
.measure tran avgvall1bl264 AVG v(l1bl264) FROM = 199ns TO =200ns
.measure tran avgvall1bl265 AVG v(l1bl265) FROM = 199ns TO =200ns
.measure tran avgvall1bl266 AVG v(l1bl266) FROM = 199ns TO =200ns
.measure tran avgvall1bl267 AVG v(l1bl267) FROM = 199ns TO =200ns
.measure tran avgvall1bl268 AVG v(l1bl268) FROM = 199ns TO =200ns
.measure tran avgvall1bl269 AVG v(l1bl269) FROM = 199ns TO =200ns
.measure tran avgvall1bl270 AVG v(l1bl270) FROM = 199ns TO =200ns
.measure tran avgvall1bl271 AVG v(l1bl271) FROM = 199ns TO =200ns
.measure tran avgvall1bl272 AVG v(l1bl272) FROM = 199ns TO =200ns
.measure tran avgvall1bl273 AVG v(l1bl273) FROM = 199ns TO =200ns
.measure tran avgvall1bl274 AVG v(l1bl274) FROM = 199ns TO =200ns
.measure tran avgvall1bl275 AVG v(l1bl275) FROM = 199ns TO =200ns
.measure tran avgvall1bl276 AVG v(l1bl276) FROM = 199ns TO =200ns
.measure tran avgvall1bl277 AVG v(l1bl277) FROM = 199ns TO =200ns
.measure tran avgvall1bl278 AVG v(l1bl278) FROM = 199ns TO =200ns
.measure tran avgvall1bl279 AVG v(l1bl279) FROM = 199ns TO =200ns
.measure tran avgvall1bl280 AVG v(l1bl280) FROM = 199ns TO =200ns
.measure tran avgvall1bl281 AVG v(l1bl281) FROM = 199ns TO =200ns
.measure tran avgvall1bl282 AVG v(l1bl282) FROM = 199ns TO =200ns
.measure tran avgvall1bl283 AVG v(l1bl283) FROM = 199ns TO =200ns
.measure tran avgvall1bl284 AVG v(l1bl284) FROM = 199ns TO =200ns
.measure tran avgvall1bl285 AVG v(l1bl285) FROM = 199ns TO =200ns
.measure tran avgvall1bl286 AVG v(l1bl286) FROM = 199ns TO =200ns
.measure tran avgvall1bl287 AVG v(l1bl287) FROM = 199ns TO =200ns
.measure tran avgvall1bl288 AVG v(l1bl288) FROM = 199ns TO =200ns
.measure tran avgvall1bl289 AVG v(l1bl289) FROM = 199ns TO =200ns
.measure tran avgvall1bl290 AVG v(l1bl290) FROM = 199ns TO =200ns
.measure tran avgvall1bl291 AVG v(l1bl291) FROM = 199ns TO =200ns
.measure tran avgvall1bl292 AVG v(l1bl292) FROM = 199ns TO =200ns
.measure tran avgvall1bl293 AVG v(l1bl293) FROM = 199ns TO =200ns
.measure tran avgvall1bl294 AVG v(l1bl294) FROM = 199ns TO =200ns
.measure tran avgvall1bl295 AVG v(l1bl295) FROM = 199ns TO =200ns
.measure tran avgvall1bl296 AVG v(l1bl296) FROM = 199ns TO =200ns
.measure tran avgvall1bl297 AVG v(l1bl297) FROM = 199ns TO =200ns
.measure tran avgvall1bl298 AVG v(l1bl298) FROM = 199ns TO =200ns
.measure tran avgvall1bl299 AVG v(l1bl299) FROM = 199ns TO =200ns
.measure tran avgvall1bl300 AVG v(l1bl300) FROM = 199ns TO =200ns
.measure tran avgvall1bl301 AVG v(l1bl301) FROM = 199ns TO =200ns
.measure tran avgvall1bl302 AVG v(l1bl302) FROM = 199ns TO =200ns
.measure tran avgvall1bl303 AVG v(l1bl303) FROM = 199ns TO =200ns
.measure tran avgvall1bl304 AVG v(l1bl304) FROM = 199ns TO =200ns
.measure tran avgvall1bl305 AVG v(l1bl305) FROM = 199ns TO =200ns
.measure tran avgvall1bl306 AVG v(l1bl306) FROM = 199ns TO =200ns
.measure tran avgvall1bl307 AVG v(l1bl307) FROM = 199ns TO =200ns
.measure tran avgvall1bl308 AVG v(l1bl308) FROM = 199ns TO =200ns
.measure tran avgvall1bl309 AVG v(l1bl309) FROM = 199ns TO =200ns
.measure tran avgvall1bl310 AVG v(l1bl310) FROM = 199ns TO =200ns
.measure tran avgvall1bl311 AVG v(l1bl311) FROM = 199ns TO =200ns
.measure tran avgvall1bl312 AVG v(l1bl312) FROM = 199ns TO =200ns
.measure tran avgvall1bl313 AVG v(l1bl313) FROM = 199ns TO =200ns
.measure tran avgvall1bl314 AVG v(l1bl314) FROM = 199ns TO =200ns
.measure tran avgvall1bl315 AVG v(l1bl315) FROM = 199ns TO =200ns
.measure tran avgvall1bl316 AVG v(l1bl316) FROM = 199ns TO =200ns
.measure tran avgvall1bl317 AVG v(l1bl317) FROM = 199ns TO =200ns
.measure tran avgvall1bl318 AVG v(l1bl318) FROM = 199ns TO =200ns
.measure tran avgvall1bl319 AVG v(l1bl319) FROM = 199ns TO =200ns
.measure tran avgvall1bl320 AVG v(l1bl320) FROM = 199ns TO =200ns
.measure tran avgvall1bl321 AVG v(l1bl321) FROM = 199ns TO =200ns
.measure tran avgvall1bl322 AVG v(l1bl322) FROM = 199ns TO =200ns
.measure tran avgvall1bl323 AVG v(l1bl323) FROM = 199ns TO =200ns
.measure tran avgvall1bl324 AVG v(l1bl324) FROM = 199ns TO =200ns
.measure tran avgvall1bl325 AVG v(l1bl325) FROM = 199ns TO =200ns
.measure tran avgvall1bl326 AVG v(l1bl326) FROM = 199ns TO =200ns
.measure tran avgvall1bl327 AVG v(l1bl327) FROM = 199ns TO =200ns
.measure tran avgvall1bl328 AVG v(l1bl328) FROM = 199ns TO =200ns
.measure tran avgvall1bl329 AVG v(l1bl329) FROM = 199ns TO =200ns
.measure tran avgvall1bl330 AVG v(l1bl330) FROM = 199ns TO =200ns
.measure tran avgvall1bl331 AVG v(l1bl331) FROM = 199ns TO =200ns
.measure tran avgvall1bl332 AVG v(l1bl332) FROM = 199ns TO =200ns
.measure tran avgvall1bl333 AVG v(l1bl333) FROM = 199ns TO =200ns
.measure tran avgvall1bl334 AVG v(l1bl334) FROM = 199ns TO =200ns
.measure tran avgvall1bl335 AVG v(l1bl335) FROM = 199ns TO =200ns
.measure tran avgvall1bl336 AVG v(l1bl336) FROM = 199ns TO =200ns
.measure tran avgvall1bl337 AVG v(l1bl337) FROM = 199ns TO =200ns
.measure tran avgvall1bl338 AVG v(l1bl338) FROM = 199ns TO =200ns
.measure tran avgvall1bl339 AVG v(l1bl339) FROM = 199ns TO =200ns
.measure tran avgvall1bl340 AVG v(l1bl340) FROM = 199ns TO =200ns
.measure tran avgvall1bl341 AVG v(l1bl341) FROM = 199ns TO =200ns
.measure tran avgvall1bl342 AVG v(l1bl342) FROM = 199ns TO =200ns
.measure tran avgvall1bl343 AVG v(l1bl343) FROM = 199ns TO =200ns
.measure tran avgvall1bl344 AVG v(l1bl344) FROM = 199ns TO =200ns
.measure tran avgvall1bl345 AVG v(l1bl345) FROM = 199ns TO =200ns
.measure tran avgvall1bl346 AVG v(l1bl346) FROM = 199ns TO =200ns
.measure tran avgvall1bl347 AVG v(l1bl347) FROM = 199ns TO =200ns
.measure tran avgvall1bl348 AVG v(l1bl348) FROM = 199ns TO =200ns
.measure tran avgvall1bl349 AVG v(l1bl349) FROM = 199ns TO =200ns
.measure tran avgvall1bl350 AVG v(l1bl350) FROM = 199ns TO =200ns
.measure tran avgvall1bl351 AVG v(l1bl351) FROM = 199ns TO =200ns
.measure tran avgvall1bl352 AVG v(l1bl352) FROM = 199ns TO =200ns
.measure tran avgvall1bl353 AVG v(l1bl353) FROM = 199ns TO =200ns
.measure tran avgvall1bl354 AVG v(l1bl354) FROM = 199ns TO =200ns
.measure tran avgvall1bl355 AVG v(l1bl355) FROM = 199ns TO =200ns
.measure tran avgvall1bl356 AVG v(l1bl356) FROM = 199ns TO =200ns
.measure tran avgvall1bl357 AVG v(l1bl357) FROM = 199ns TO =200ns
.measure tran avgvall1bl358 AVG v(l1bl358) FROM = 199ns TO =200ns
.measure tran avgvall1bl359 AVG v(l1bl359) FROM = 199ns TO =200ns
.measure tran avgvall1bl360 AVG v(l1bl360) FROM = 199ns TO =200ns
.measure tran avgvall1bl361 AVG v(l1bl361) FROM = 199ns TO =200ns
.measure tran avgvall1bl362 AVG v(l1bl362) FROM = 199ns TO =200ns
.measure tran avgvall1bl363 AVG v(l1bl363) FROM = 199ns TO =200ns
.measure tran avgvall1bl364 AVG v(l1bl364) FROM = 199ns TO =200ns
.measure tran avgvall1bl365 AVG v(l1bl365) FROM = 199ns TO =200ns
.measure tran avgvall1bl366 AVG v(l1bl366) FROM = 199ns TO =200ns
.measure tran avgvall1bl367 AVG v(l1bl367) FROM = 199ns TO =200ns
.measure tran avgvall1bl368 AVG v(l1bl368) FROM = 199ns TO =200ns
.measure tran avgvall1bl369 AVG v(l1bl369) FROM = 199ns TO =200ns
.measure tran avgvall1bl370 AVG v(l1bl370) FROM = 199ns TO =200ns
.measure tran avgvall1bl371 AVG v(l1bl371) FROM = 199ns TO =200ns
.measure tran avgvall1bl372 AVG v(l1bl372) FROM = 199ns TO =200ns
.measure tran avgvall1bl373 AVG v(l1bl373) FROM = 199ns TO =200ns
.measure tran avgvall1bl374 AVG v(l1bl374) FROM = 199ns TO =200ns
.measure tran avgvall1bl375 AVG v(l1bl375) FROM = 199ns TO =200ns
.measure tran avgvall1bl376 AVG v(l1bl376) FROM = 199ns TO =200ns
.measure tran avgvall1bl377 AVG v(l1bl377) FROM = 199ns TO =200ns
.measure tran avgvall1bl378 AVG v(l1bl378) FROM = 199ns TO =200ns
.measure tran avgvall1bl379 AVG v(l1bl379) FROM = 199ns TO =200ns
.measure tran avgvall1bl380 AVG v(l1bl380) FROM = 199ns TO =200ns
.measure tran avgvall1bl381 AVG v(l1bl381) FROM = 199ns TO =200ns
.measure tran avgvall1bl382 AVG v(l1bl382) FROM = 199ns TO =200ns
.measure tran avgvall1bl383 AVG v(l1bl383) FROM = 199ns TO =200ns
.measure tran avgvall1bl384 AVG v(l1bl384) FROM = 199ns TO =200ns
.measure tran avgvall1bl385 AVG v(l1bl385) FROM = 199ns TO =200ns
.measure tran avgvall1bl386 AVG v(l1bl386) FROM = 199ns TO =200ns
.measure tran avgvall1bl387 AVG v(l1bl387) FROM = 199ns TO =200ns
.measure tran avgvall1bl388 AVG v(l1bl388) FROM = 199ns TO =200ns
.measure tran avgvall1bl389 AVG v(l1bl389) FROM = 199ns TO =200ns
.measure tran avgvall1bl390 AVG v(l1bl390) FROM = 199ns TO =200ns
.measure tran avgvall1bl391 AVG v(l1bl391) FROM = 199ns TO =200ns
.measure tran avgvall1bl392 AVG v(l1bl392) FROM = 199ns TO =200ns
.measure tran avgvall1bl393 AVG v(l1bl393) FROM = 199ns TO =200ns
.measure tran avgvall1bl394 AVG v(l1bl394) FROM = 199ns TO =200ns
.measure tran avgvall1bl395 AVG v(l1bl395) FROM = 199ns TO =200ns
.measure tran avgvall1bl396 AVG v(l1bl396) FROM = 199ns TO =200ns
.measure tran avgvall1bl397 AVG v(l1bl397) FROM = 199ns TO =200ns
.measure tran avgvall1bl398 AVG v(l1bl398) FROM = 199ns TO =200ns
.measure tran avgvall1bl399 AVG v(l1bl399) FROM = 199ns TO =200ns
.measure tran avgvall1bl400 AVG v(l1bl400) FROM = 199ns TO =200ns
.measure tran avgvall1bl401 AVG v(l1bl401) FROM = 199ns TO =200ns
.measure tran avgvall1bl402 AVG v(l1bl402) FROM = 199ns TO =200ns
.measure tran avgvall1bl403 AVG v(l1bl403) FROM = 199ns TO =200ns
.measure tran avgvall1bl404 AVG v(l1bl404) FROM = 199ns TO =200ns
.measure tran avgvall1bl405 AVG v(l1bl405) FROM = 199ns TO =200ns
.measure tran avgvall1bl406 AVG v(l1bl406) FROM = 199ns TO =200ns
.measure tran avgvall1bl407 AVG v(l1bl407) FROM = 199ns TO =200ns
.measure tran avgvall1bl408 AVG v(l1bl408) FROM = 199ns TO =200ns
.measure tran avgvall1bl409 AVG v(l1bl409) FROM = 199ns TO =200ns
.measure tran avgvall1bl410 AVG v(l1bl410) FROM = 199ns TO =200ns
.measure tran avgvall1bl411 AVG v(l1bl411) FROM = 199ns TO =200ns
.measure tran avgvall1bl412 AVG v(l1bl412) FROM = 199ns TO =200ns
.measure tran avgvall1bl413 AVG v(l1bl413) FROM = 199ns TO =200ns
.measure tran avgvall1bl414 AVG v(l1bl414) FROM = 199ns TO =200ns
.measure tran avgvall1bl415 AVG v(l1bl415) FROM = 199ns TO =200ns
.measure tran avgvall1bl416 AVG v(l1bl416) FROM = 199ns TO =200ns
.measure tran avgvall1bl417 AVG v(l1bl417) FROM = 199ns TO =200ns
.measure tran avgvall1bl418 AVG v(l1bl418) FROM = 199ns TO =200ns
.measure tran avgvall1bl419 AVG v(l1bl419) FROM = 199ns TO =200ns
.measure tran avgvall1bl420 AVG v(l1bl420) FROM = 199ns TO =200ns
.measure tran avgvall1bl421 AVG v(l1bl421) FROM = 199ns TO =200ns
.measure tran avgvall1bl422 AVG v(l1bl422) FROM = 199ns TO =200ns
.measure tran avgvall1bl423 AVG v(l1bl423) FROM = 199ns TO =200ns
.measure tran avgvall1bl424 AVG v(l1bl424) FROM = 199ns TO =200ns
.measure tran avgvall1bl425 AVG v(l1bl425) FROM = 199ns TO =200ns
.measure tran avgvall1bl426 AVG v(l1bl426) FROM = 199ns TO =200ns
.measure tran avgvall1bl427 AVG v(l1bl427) FROM = 199ns TO =200ns
.measure tran avgvall1bl428 AVG v(l1bl428) FROM = 199ns TO =200ns
.measure tran avgvall1bl429 AVG v(l1bl429) FROM = 199ns TO =200ns
.measure tran avgvall1bl430 AVG v(l1bl430) FROM = 199ns TO =200ns
.measure tran avgvall1bl431 AVG v(l1bl431) FROM = 199ns TO =200ns
.measure tran avgvall1bl432 AVG v(l1bl432) FROM = 199ns TO =200ns
.measure tran avgvall1bl433 AVG v(l1bl433) FROM = 199ns TO =200ns
.measure tran avgvall1bl434 AVG v(l1bl434) FROM = 199ns TO =200ns
.measure tran avgvall1bl435 AVG v(l1bl435) FROM = 199ns TO =200ns
.measure tran avgvall1bl436 AVG v(l1bl436) FROM = 199ns TO =200ns
.measure tran avgvall1bl437 AVG v(l1bl437) FROM = 199ns TO =200ns
.measure tran avgvall1bl438 AVG v(l1bl438) FROM = 199ns TO =200ns
.measure tran avgvall1bl439 AVG v(l1bl439) FROM = 199ns TO =200ns
.measure tran avgvall1bl440 AVG v(l1bl440) FROM = 199ns TO =200ns
.measure tran avgvall1bl441 AVG v(l1bl441) FROM = 199ns TO =200ns
.measure tran avgvall1bl442 AVG v(l1bl442) FROM = 199ns TO =200ns
.measure tran avgvall1bl443 AVG v(l1bl443) FROM = 199ns TO =200ns
.measure tran avgvall1bl444 AVG v(l1bl444) FROM = 199ns TO =200ns
.measure tran avgvall1bl445 AVG v(l1bl445) FROM = 199ns TO =200ns
.measure tran avgvall1bl446 AVG v(l1bl446) FROM = 199ns TO =200ns
.measure tran avgvall1bl447 AVG v(l1bl447) FROM = 199ns TO =200ns
.measure tran avgvall1bl448 AVG v(l1bl448) FROM = 199ns TO =200ns
.measure tran avgvall1bl449 AVG v(l1bl449) FROM = 199ns TO =200ns
.measure tran avgvall1bl450 AVG v(l1bl450) FROM = 199ns TO =200ns
.measure tran avgvall1bl451 AVG v(l1bl451) FROM = 199ns TO =200ns
.measure tran avgvall1bl452 AVG v(l1bl452) FROM = 199ns TO =200ns
.measure tran avgvall1bl453 AVG v(l1bl453) FROM = 199ns TO =200ns
.measure tran avgvall1bl454 AVG v(l1bl454) FROM = 199ns TO =200ns
.measure tran avgvall1bl455 AVG v(l1bl455) FROM = 199ns TO =200ns
.measure tran avgvall1bl456 AVG v(l1bl456) FROM = 199ns TO =200ns
.measure tran avgvall1bl457 AVG v(l1bl457) FROM = 199ns TO =200ns
.measure tran avgvall1bl458 AVG v(l1bl458) FROM = 199ns TO =200ns
.measure tran avgvall1bl459 AVG v(l1bl459) FROM = 199ns TO =200ns
.measure tran avgvall1bl460 AVG v(l1bl460) FROM = 199ns TO =200ns
.measure tran avgvall1bl461 AVG v(l1bl461) FROM = 199ns TO =200ns
.measure tran avgvall1bl462 AVG v(l1bl462) FROM = 199ns TO =200ns
.measure tran avgvall1bl463 AVG v(l1bl463) FROM = 199ns TO =200ns
.measure tran avgvall1bl464 AVG v(l1bl464) FROM = 199ns TO =200ns
.measure tran avgvall1bl465 AVG v(l1bl465) FROM = 199ns TO =200ns
.measure tran avgvall1bl466 AVG v(l1bl466) FROM = 199ns TO =200ns
.measure tran avgvall1bl467 AVG v(l1bl467) FROM = 199ns TO =200ns
.measure tran avgvall1bl468 AVG v(l1bl468) FROM = 199ns TO =200ns
.measure tran avgvall1bl469 AVG v(l1bl469) FROM = 199ns TO =200ns
.measure tran avgvall1bl470 AVG v(l1bl470) FROM = 199ns TO =200ns
.measure tran avgvall1bl471 AVG v(l1bl471) FROM = 199ns TO =200ns
.measure tran avgvall1bl472 AVG v(l1bl472) FROM = 199ns TO =200ns
.measure tran avgvall1bl473 AVG v(l1bl473) FROM = 199ns TO =200ns
.measure tran avgvall1bl474 AVG v(l1bl474) FROM = 199ns TO =200ns
.measure tran avgvall1bl475 AVG v(l1bl475) FROM = 199ns TO =200ns
.measure tran avgvall1bl476 AVG v(l1bl476) FROM = 199ns TO =200ns
.measure tran avgvall1bl477 AVG v(l1bl477) FROM = 199ns TO =200ns
.measure tran avgvall1bl478 AVG v(l1bl478) FROM = 199ns TO =200ns
.measure tran avgvall1bl479 AVG v(l1bl479) FROM = 199ns TO =200ns
.measure tran avgvall1bl480 AVG v(l1bl480) FROM = 199ns TO =200ns
.measure tran avgvall1bl481 AVG v(l1bl481) FROM = 199ns TO =200ns
.measure tran avgvall1bl482 AVG v(l1bl482) FROM = 199ns TO =200ns
.measure tran avgvall1bl483 AVG v(l1bl483) FROM = 199ns TO =200ns
.measure tran avgvall1bl484 AVG v(l1bl484) FROM = 199ns TO =200ns
.measure tran avgvall1bl485 AVG v(l1bl485) FROM = 199ns TO =200ns
.measure tran avgvall1bl486 AVG v(l1bl486) FROM = 199ns TO =200ns
.measure tran avgvall1bl487 AVG v(l1bl487) FROM = 199ns TO =200ns
.measure tran avgvall1bl488 AVG v(l1bl488) FROM = 199ns TO =200ns
.measure tran avgvall1bl489 AVG v(l1bl489) FROM = 199ns TO =200ns
.measure tran avgvall1bl490 AVG v(l1bl490) FROM = 199ns TO =200ns
.measure tran avgvall1bl491 AVG v(l1bl491) FROM = 199ns TO =200ns
.measure tran avgvall1bl492 AVG v(l1bl492) FROM = 199ns TO =200ns
.measure tran avgvall1bl493 AVG v(l1bl493) FROM = 199ns TO =200ns
.measure tran avgvall1bl494 AVG v(l1bl494) FROM = 199ns TO =200ns
.measure tran avgvall1bl495 AVG v(l1bl495) FROM = 199ns TO =200ns
.measure tran avgvall1bl496 AVG v(l1bl496) FROM = 199ns TO =200ns
.measure tran avgvall1bl497 AVG v(l1bl497) FROM = 199ns TO =200ns
.measure tran avgvall1bl498 AVG v(l1bl498) FROM = 199ns TO =200ns
.measure tran avgvall1bl499 AVG v(l1bl499) FROM = 199ns TO =200ns
.measure tran avgvall1bl500 AVG v(l1bl500) FROM = 199ns TO =200ns
.measure tran avgvall1bl501 AVG v(l1bl501) FROM = 199ns TO =200ns
.measure tran avgvall1bl502 AVG v(l1bl502) FROM = 199ns TO =200ns
.measure tran avgvall1bl503 AVG v(l1bl503) FROM = 199ns TO =200ns
.measure tran avgvall1bl504 AVG v(l1bl504) FROM = 199ns TO =200ns
.measure tran avgvall1bl505 AVG v(l1bl505) FROM = 199ns TO =200ns
.measure tran avgvall1bl506 AVG v(l1bl506) FROM = 199ns TO =200ns
.measure tran avgvall1bl507 AVG v(l1bl507) FROM = 199ns TO =200ns
.measure tran avgvall1bl508 AVG v(l1bl508) FROM = 199ns TO =200ns
.measure tran avgvall1bl509 AVG v(l1bl509) FROM = 199ns TO =200ns
.measure tran avgvall1bl510 AVG v(l1bl510) FROM = 199ns TO =200ns
.measure tran avgvall1bl511 AVG v(l1bl511) FROM = 199ns TO =200ns

.measure tran avgvall2bl0 AVG v(l2bl0) FROM = 199ns TO =200ns
.measure tran avgvall2bl1 AVG v(l2bl1) FROM = 199ns TO =200ns
.measure tran avgvall2bl2 AVG v(l2bl2) FROM = 199ns TO =200ns
.measure tran avgvall2bl3 AVG v(l2bl3) FROM = 199ns TO =200ns
.measure tran avgvall2bl4 AVG v(l2bl4) FROM = 199ns TO =200ns
.measure tran avgvall2bl5 AVG v(l2bl5) FROM = 199ns TO =200ns
.measure tran avgvall2bl6 AVG v(l2bl6) FROM = 199ns TO =200ns
.measure tran avgvall2bl7 AVG v(l2bl7) FROM = 199ns TO =200ns
.measure tran avgvall2bl8 AVG v(l2bl8) FROM = 199ns TO =200ns
.measure tran avgvall2bl9 AVG v(l2bl9) FROM = 199ns TO =200ns
.measure tran avgvall2bl10 AVG v(l2bl10) FROM = 199ns TO =200ns
.measure tran avgvall2bl11 AVG v(l2bl11) FROM = 199ns TO =200ns
.measure tran avgvall2bl12 AVG v(l2bl12) FROM = 199ns TO =200ns
.measure tran avgvall2bl13 AVG v(l2bl13) FROM = 199ns TO =200ns
.measure tran avgvall2bl14 AVG v(l2bl14) FROM = 199ns TO =200ns
.measure tran avgvall2bl15 AVG v(l2bl15) FROM = 199ns TO =200ns
.measure tran avgvall2bl16 AVG v(l2bl16) FROM = 199ns TO =200ns
.measure tran avgvall2bl17 AVG v(l2bl17) FROM = 199ns TO =200ns
.measure tran avgvall2bl18 AVG v(l2bl18) FROM = 199ns TO =200ns
.measure tran avgvall2bl19 AVG v(l2bl19) FROM = 199ns TO =200ns
.measure tran avgvall2bl20 AVG v(l2bl20) FROM = 199ns TO =200ns
.measure tran avgvall2bl21 AVG v(l2bl21) FROM = 199ns TO =200ns
.measure tran avgvall2bl22 AVG v(l2bl22) FROM = 199ns TO =200ns
.measure tran avgvall2bl23 AVG v(l2bl23) FROM = 199ns TO =200ns
.measure tran avgvall2bl24 AVG v(l2bl24) FROM = 199ns TO =200ns
.measure tran avgvall2bl25 AVG v(l2bl25) FROM = 199ns TO =200ns
.measure tran avgvall2bl26 AVG v(l2bl26) FROM = 199ns TO =200ns
.measure tran avgvall2bl27 AVG v(l2bl27) FROM = 199ns TO =200ns
.measure tran avgvall2bl28 AVG v(l2bl28) FROM = 199ns TO =200ns
.measure tran avgvall2bl29 AVG v(l2bl29) FROM = 199ns TO =200ns
.measure tran avgvall2bl30 AVG v(l2bl30) FROM = 199ns TO =200ns
.measure tran avgvall2bl31 AVG v(l2bl31) FROM = 199ns TO =200ns
.measure tran avgvall2bl32 AVG v(l2bl32) FROM = 199ns TO =200ns
.measure tran avgvall2bl33 AVG v(l2bl33) FROM = 199ns TO =200ns
.measure tran avgvall2bl34 AVG v(l2bl34) FROM = 199ns TO =200ns
.measure tran avgvall2bl35 AVG v(l2bl35) FROM = 199ns TO =200ns
.measure tran avgvall2bl36 AVG v(l2bl36) FROM = 199ns TO =200ns
.measure tran avgvall2bl37 AVG v(l2bl37) FROM = 199ns TO =200ns
.measure tran avgvall2bl38 AVG v(l2bl38) FROM = 199ns TO =200ns
.measure tran avgvall2bl39 AVG v(l2bl39) FROM = 199ns TO =200ns
.measure tran avgvall2bl40 AVG v(l2bl40) FROM = 199ns TO =200ns
.measure tran avgvall2bl41 AVG v(l2bl41) FROM = 199ns TO =200ns
.measure tran avgvall2bl42 AVG v(l2bl42) FROM = 199ns TO =200ns
.measure tran avgvall2bl43 AVG v(l2bl43) FROM = 199ns TO =200ns
.measure tran avgvall2bl44 AVG v(l2bl44) FROM = 199ns TO =200ns
.measure tran avgvall2bl45 AVG v(l2bl45) FROM = 199ns TO =200ns
.measure tran avgvall2bl46 AVG v(l2bl46) FROM = 199ns TO =200ns
.measure tran avgvall2bl47 AVG v(l2bl47) FROM = 199ns TO =200ns
.measure tran avgvall2bl48 AVG v(l2bl48) FROM = 199ns TO =200ns
.measure tran avgvall2bl49 AVG v(l2bl49) FROM = 199ns TO =200ns
.measure tran avgvall2bl50 AVG v(l2bl50) FROM = 199ns TO =200ns
.measure tran avgvall2bl51 AVG v(l2bl51) FROM = 199ns TO =200ns
.measure tran avgvall2bl52 AVG v(l2bl52) FROM = 199ns TO =200ns
.measure tran avgvall2bl53 AVG v(l2bl53) FROM = 199ns TO =200ns
.measure tran avgvall2bl54 AVG v(l2bl54) FROM = 199ns TO =200ns
.measure tran avgvall2bl55 AVG v(l2bl55) FROM = 199ns TO =200ns
.measure tran avgvall2bl56 AVG v(l2bl56) FROM = 199ns TO =200ns
.measure tran avgvall2bl57 AVG v(l2bl57) FROM = 199ns TO =200ns
.measure tran avgvall2bl58 AVG v(l2bl58) FROM = 199ns TO =200ns
.measure tran avgvall2bl59 AVG v(l2bl59) FROM = 199ns TO =200ns
.measure tran avgvall2bl60 AVG v(l2bl60) FROM = 199ns TO =200ns
.measure tran avgvall2bl61 AVG v(l2bl61) FROM = 199ns TO =200ns
.measure tran avgvall2bl62 AVG v(l2bl62) FROM = 199ns TO =200ns
.measure tran avgvall2bl63 AVG v(l2bl63) FROM = 199ns TO =200ns
.measure tran avgvall2bl64 AVG v(l2bl64) FROM = 199ns TO =200ns
.measure tran avgvall2bl65 AVG v(l2bl65) FROM = 199ns TO =200ns
.measure tran avgvall2bl66 AVG v(l2bl66) FROM = 199ns TO =200ns
.measure tran avgvall2bl67 AVG v(l2bl67) FROM = 199ns TO =200ns
.measure tran avgvall2bl68 AVG v(l2bl68) FROM = 199ns TO =200ns
.measure tran avgvall2bl69 AVG v(l2bl69) FROM = 199ns TO =200ns
.measure tran avgvall2bl70 AVG v(l2bl70) FROM = 199ns TO =200ns
.measure tran avgvall2bl71 AVG v(l2bl71) FROM = 199ns TO =200ns
.measure tran avgvall2bl72 AVG v(l2bl72) FROM = 199ns TO =200ns
.measure tran avgvall2bl73 AVG v(l2bl73) FROM = 199ns TO =200ns
.measure tran avgvall2bl74 AVG v(l2bl74) FROM = 199ns TO =200ns
.measure tran avgvall2bl75 AVG v(l2bl75) FROM = 199ns TO =200ns
.measure tran avgvall2bl76 AVG v(l2bl76) FROM = 199ns TO =200ns
.measure tran avgvall2bl77 AVG v(l2bl77) FROM = 199ns TO =200ns
.measure tran avgvall2bl78 AVG v(l2bl78) FROM = 199ns TO =200ns
.measure tran avgvall2bl79 AVG v(l2bl79) FROM = 199ns TO =200ns
.measure tran avgvall2bl80 AVG v(l2bl80) FROM = 199ns TO =200ns
.measure tran avgvall2bl81 AVG v(l2bl81) FROM = 199ns TO =200ns
.measure tran avgvall2bl82 AVG v(l2bl82) FROM = 199ns TO =200ns
.measure tran avgvall2bl83 AVG v(l2bl83) FROM = 199ns TO =200ns
.measure tran avgvall2bl84 AVG v(l2bl84) FROM = 199ns TO =200ns
.measure tran avgvall2bl85 AVG v(l2bl85) FROM = 199ns TO =200ns
.measure tran avgvall2bl86 AVG v(l2bl86) FROM = 199ns TO =200ns
.measure tran avgvall2bl87 AVG v(l2bl87) FROM = 199ns TO =200ns
.measure tran avgvall2bl88 AVG v(l2bl88) FROM = 199ns TO =200ns
.measure tran avgvall2bl89 AVG v(l2bl89) FROM = 199ns TO =200ns
.measure tran avgvall2bl90 AVG v(l2bl90) FROM = 199ns TO =200ns
.measure tran avgvall2bl91 AVG v(l2bl91) FROM = 199ns TO =200ns
.measure tran avgvall2bl92 AVG v(l2bl92) FROM = 199ns TO =200ns
.measure tran avgvall2bl93 AVG v(l2bl93) FROM = 199ns TO =200ns
.measure tran avgvall2bl94 AVG v(l2bl94) FROM = 199ns TO =200ns
.measure tran avgvall2bl95 AVG v(l2bl95) FROM = 199ns TO =200ns
.measure tran avgvall2bl96 AVG v(l2bl96) FROM = 199ns TO =200ns
.measure tran avgvall2bl97 AVG v(l2bl97) FROM = 199ns TO =200ns
.measure tran avgvall2bl98 AVG v(l2bl98) FROM = 199ns TO =200ns
.measure tran avgvall2bl99 AVG v(l2bl99) FROM = 199ns TO =200ns
.measure tran avgvall2bl100 AVG v(l2bl100) FROM = 199ns TO =200ns
.measure tran avgvall2bl101 AVG v(l2bl101) FROM = 199ns TO =200ns
.measure tran avgvall2bl102 AVG v(l2bl102) FROM = 199ns TO =200ns
.measure tran avgvall2bl103 AVG v(l2bl103) FROM = 199ns TO =200ns
.measure tran avgvall2bl104 AVG v(l2bl104) FROM = 199ns TO =200ns
.measure tran avgvall2bl105 AVG v(l2bl105) FROM = 199ns TO =200ns
.measure tran avgvall2bl106 AVG v(l2bl106) FROM = 199ns TO =200ns
.measure tran avgvall2bl107 AVG v(l2bl107) FROM = 199ns TO =200ns
.measure tran avgvall2bl108 AVG v(l2bl108) FROM = 199ns TO =200ns
.measure tran avgvall2bl109 AVG v(l2bl109) FROM = 199ns TO =200ns
.measure tran avgvall2bl110 AVG v(l2bl110) FROM = 199ns TO =200ns
.measure tran avgvall2bl111 AVG v(l2bl111) FROM = 199ns TO =200ns
.measure tran avgvall2bl112 AVG v(l2bl112) FROM = 199ns TO =200ns
.measure tran avgvall2bl113 AVG v(l2bl113) FROM = 199ns TO =200ns
.measure tran avgvall2bl114 AVG v(l2bl114) FROM = 199ns TO =200ns
.measure tran avgvall2bl115 AVG v(l2bl115) FROM = 199ns TO =200ns
.measure tran avgvall2bl116 AVG v(l2bl116) FROM = 199ns TO =200ns
.measure tran avgvall2bl117 AVG v(l2bl117) FROM = 199ns TO =200ns
.measure tran avgvall2bl118 AVG v(l2bl118) FROM = 199ns TO =200ns
.measure tran avgvall2bl119 AVG v(l2bl119) FROM = 199ns TO =200ns
.measure tran avgvall2bl120 AVG v(l2bl120) FROM = 199ns TO =200ns
.measure tran avgvall2bl121 AVG v(l2bl121) FROM = 199ns TO =200ns
.measure tran avgvall2bl122 AVG v(l2bl122) FROM = 199ns TO =200ns
.measure tran avgvall2bl123 AVG v(l2bl123) FROM = 199ns TO =200ns
.measure tran avgvall2bl124 AVG v(l2bl124) FROM = 199ns TO =200ns
.measure tran avgvall2bl125 AVG v(l2bl125) FROM = 199ns TO =200ns
.measure tran avgvall2bl126 AVG v(l2bl126) FROM = 199ns TO =200ns
.measure tran avgvall2bl127 AVG v(l2bl127) FROM = 199ns TO =200ns
.measure tran avgvall2bl128 AVG v(l2bl128) FROM = 199ns TO =200ns
.measure tran avgvall2bl129 AVG v(l2bl129) FROM = 199ns TO =200ns
.measure tran avgvall2bl130 AVG v(l2bl130) FROM = 199ns TO =200ns
.measure tran avgvall2bl131 AVG v(l2bl131) FROM = 199ns TO =200ns
.measure tran avgvall2bl132 AVG v(l2bl132) FROM = 199ns TO =200ns
.measure tran avgvall2bl133 AVG v(l2bl133) FROM = 199ns TO =200ns
.measure tran avgvall2bl134 AVG v(l2bl134) FROM = 199ns TO =200ns
.measure tran avgvall2bl135 AVG v(l2bl135) FROM = 199ns TO =200ns
.measure tran avgvall2bl136 AVG v(l2bl136) FROM = 199ns TO =200ns
.measure tran avgvall2bl137 AVG v(l2bl137) FROM = 199ns TO =200ns
.measure tran avgvall2bl138 AVG v(l2bl138) FROM = 199ns TO =200ns
.measure tran avgvall2bl139 AVG v(l2bl139) FROM = 199ns TO =200ns
.measure tran avgvall2bl140 AVG v(l2bl140) FROM = 199ns TO =200ns
.measure tran avgvall2bl141 AVG v(l2bl141) FROM = 199ns TO =200ns
.measure tran avgvall2bl142 AVG v(l2bl142) FROM = 199ns TO =200ns
.measure tran avgvall2bl143 AVG v(l2bl143) FROM = 199ns TO =200ns
.measure tran avgvall2bl144 AVG v(l2bl144) FROM = 199ns TO =200ns
.measure tran avgvall2bl145 AVG v(l2bl145) FROM = 199ns TO =200ns
.measure tran avgvall2bl146 AVG v(l2bl146) FROM = 199ns TO =200ns
.measure tran avgvall2bl147 AVG v(l2bl147) FROM = 199ns TO =200ns
.measure tran avgvall2bl148 AVG v(l2bl148) FROM = 199ns TO =200ns
.measure tran avgvall2bl149 AVG v(l2bl149) FROM = 199ns TO =200ns
.measure tran avgvall2bl150 AVG v(l2bl150) FROM = 199ns TO =200ns
.measure tran avgvall2bl151 AVG v(l2bl151) FROM = 199ns TO =200ns
.measure tran avgvall2bl152 AVG v(l2bl152) FROM = 199ns TO =200ns
.measure tran avgvall2bl153 AVG v(l2bl153) FROM = 199ns TO =200ns
.measure tran avgvall2bl154 AVG v(l2bl154) FROM = 199ns TO =200ns
.measure tran avgvall2bl155 AVG v(l2bl155) FROM = 199ns TO =200ns
.measure tran avgvall2bl156 AVG v(l2bl156) FROM = 199ns TO =200ns
.measure tran avgvall2bl157 AVG v(l2bl157) FROM = 199ns TO =200ns
.measure tran avgvall2bl158 AVG v(l2bl158) FROM = 199ns TO =200ns
.measure tran avgvall2bl159 AVG v(l2bl159) FROM = 199ns TO =200ns
.measure tran avgvall2bl160 AVG v(l2bl160) FROM = 199ns TO =200ns
.measure tran avgvall2bl161 AVG v(l2bl161) FROM = 199ns TO =200ns
.measure tran avgvall2bl162 AVG v(l2bl162) FROM = 199ns TO =200ns
.measure tran avgvall2bl163 AVG v(l2bl163) FROM = 199ns TO =200ns
.measure tran avgvall2bl164 AVG v(l2bl164) FROM = 199ns TO =200ns
.measure tran avgvall2bl165 AVG v(l2bl165) FROM = 199ns TO =200ns
.measure tran avgvall2bl166 AVG v(l2bl166) FROM = 199ns TO =200ns
.measure tran avgvall2bl167 AVG v(l2bl167) FROM = 199ns TO =200ns
.measure tran avgvall2bl168 AVG v(l2bl168) FROM = 199ns TO =200ns
.measure tran avgvall2bl169 AVG v(l2bl169) FROM = 199ns TO =200ns
.measure tran avgvall2bl170 AVG v(l2bl170) FROM = 199ns TO =200ns
.measure tran avgvall2bl171 AVG v(l2bl171) FROM = 199ns TO =200ns
.measure tran avgvall2bl172 AVG v(l2bl172) FROM = 199ns TO =200ns
.measure tran avgvall2bl173 AVG v(l2bl173) FROM = 199ns TO =200ns
.measure tran avgvall2bl174 AVG v(l2bl174) FROM = 199ns TO =200ns
.measure tran avgvall2bl175 AVG v(l2bl175) FROM = 199ns TO =200ns
.measure tran avgvall2bl176 AVG v(l2bl176) FROM = 199ns TO =200ns
.measure tran avgvall2bl177 AVG v(l2bl177) FROM = 199ns TO =200ns
.measure tran avgvall2bl178 AVG v(l2bl178) FROM = 199ns TO =200ns
.measure tran avgvall2bl179 AVG v(l2bl179) FROM = 199ns TO =200ns
.measure tran avgvall2bl180 AVG v(l2bl180) FROM = 199ns TO =200ns
.measure tran avgvall2bl181 AVG v(l2bl181) FROM = 199ns TO =200ns
.measure tran avgvall2bl182 AVG v(l2bl182) FROM = 199ns TO =200ns
.measure tran avgvall2bl183 AVG v(l2bl183) FROM = 199ns TO =200ns
.measure tran avgvall2bl184 AVG v(l2bl184) FROM = 199ns TO =200ns
.measure tran avgvall2bl185 AVG v(l2bl185) FROM = 199ns TO =200ns
.measure tran avgvall2bl186 AVG v(l2bl186) FROM = 199ns TO =200ns
.measure tran avgvall2bl187 AVG v(l2bl187) FROM = 199ns TO =200ns
.measure tran avgvall2bl188 AVG v(l2bl188) FROM = 199ns TO =200ns
.measure tran avgvall2bl189 AVG v(l2bl189) FROM = 199ns TO =200ns
.measure tran avgvall2bl190 AVG v(l2bl190) FROM = 199ns TO =200ns
.measure tran avgvall2bl191 AVG v(l2bl191) FROM = 199ns TO =200ns
.measure tran avgvall2bl192 AVG v(l2bl192) FROM = 199ns TO =200ns
.measure tran avgvall2bl193 AVG v(l2bl193) FROM = 199ns TO =200ns
.measure tran avgvall2bl194 AVG v(l2bl194) FROM = 199ns TO =200ns
.measure tran avgvall2bl195 AVG v(l2bl195) FROM = 199ns TO =200ns
.measure tran avgvall2bl196 AVG v(l2bl196) FROM = 199ns TO =200ns
.measure tran avgvall2bl197 AVG v(l2bl197) FROM = 199ns TO =200ns
.measure tran avgvall2bl198 AVG v(l2bl198) FROM = 199ns TO =200ns
.measure tran avgvall2bl199 AVG v(l2bl199) FROM = 199ns TO =200ns
.measure tran avgvall2bl200 AVG v(l2bl200) FROM = 199ns TO =200ns
.measure tran avgvall2bl201 AVG v(l2bl201) FROM = 199ns TO =200ns
.measure tran avgvall2bl202 AVG v(l2bl202) FROM = 199ns TO =200ns
.measure tran avgvall2bl203 AVG v(l2bl203) FROM = 199ns TO =200ns
.measure tran avgvall2bl204 AVG v(l2bl204) FROM = 199ns TO =200ns
.measure tran avgvall2bl205 AVG v(l2bl205) FROM = 199ns TO =200ns
.measure tran avgvall2bl206 AVG v(l2bl206) FROM = 199ns TO =200ns
.measure tran avgvall2bl207 AVG v(l2bl207) FROM = 199ns TO =200ns
.measure tran avgvall2bl208 AVG v(l2bl208) FROM = 199ns TO =200ns
.measure tran avgvall2bl209 AVG v(l2bl209) FROM = 199ns TO =200ns
.measure tran avgvall2bl210 AVG v(l2bl210) FROM = 199ns TO =200ns
.measure tran avgvall2bl211 AVG v(l2bl211) FROM = 199ns TO =200ns
.measure tran avgvall2bl212 AVG v(l2bl212) FROM = 199ns TO =200ns
.measure tran avgvall2bl213 AVG v(l2bl213) FROM = 199ns TO =200ns
.measure tran avgvall2bl214 AVG v(l2bl214) FROM = 199ns TO =200ns
.measure tran avgvall2bl215 AVG v(l2bl215) FROM = 199ns TO =200ns
.measure tran avgvall2bl216 AVG v(l2bl216) FROM = 199ns TO =200ns
.measure tran avgvall2bl217 AVG v(l2bl217) FROM = 199ns TO =200ns
.measure tran avgvall2bl218 AVG v(l2bl218) FROM = 199ns TO =200ns
.measure tran avgvall2bl219 AVG v(l2bl219) FROM = 199ns TO =200ns
.measure tran avgvall2bl220 AVG v(l2bl220) FROM = 199ns TO =200ns
.measure tran avgvall2bl221 AVG v(l2bl221) FROM = 199ns TO =200ns
.measure tran avgvall2bl222 AVG v(l2bl222) FROM = 199ns TO =200ns
.measure tran avgvall2bl223 AVG v(l2bl223) FROM = 199ns TO =200ns
.measure tran avgvall2bl224 AVG v(l2bl224) FROM = 199ns TO =200ns
.measure tran avgvall2bl225 AVG v(l2bl225) FROM = 199ns TO =200ns
.measure tran avgvall2bl226 AVG v(l2bl226) FROM = 199ns TO =200ns
.measure tran avgvall2bl227 AVG v(l2bl227) FROM = 199ns TO =200ns
.measure tran avgvall2bl228 AVG v(l2bl228) FROM = 199ns TO =200ns
.measure tran avgvall2bl229 AVG v(l2bl229) FROM = 199ns TO =200ns
.measure tran avgvall2bl230 AVG v(l2bl230) FROM = 199ns TO =200ns
.measure tran avgvall2bl231 AVG v(l2bl231) FROM = 199ns TO =200ns
.measure tran avgvall2bl232 AVG v(l2bl232) FROM = 199ns TO =200ns
.measure tran avgvall2bl233 AVG v(l2bl233) FROM = 199ns TO =200ns
.measure tran avgvall2bl234 AVG v(l2bl234) FROM = 199ns TO =200ns
.measure tran avgvall2bl235 AVG v(l2bl235) FROM = 199ns TO =200ns
.measure tran avgvall2bl236 AVG v(l2bl236) FROM = 199ns TO =200ns
.measure tran avgvall2bl237 AVG v(l2bl237) FROM = 199ns TO =200ns
.measure tran avgvall2bl238 AVG v(l2bl238) FROM = 199ns TO =200ns
.measure tran avgvall2bl239 AVG v(l2bl239) FROM = 199ns TO =200ns
.measure tran avgvall2bl240 AVG v(l2bl240) FROM = 199ns TO =200ns
.measure tran avgvall2bl241 AVG v(l2bl241) FROM = 199ns TO =200ns
.measure tran avgvall2bl242 AVG v(l2bl242) FROM = 199ns TO =200ns
.measure tran avgvall2bl243 AVG v(l2bl243) FROM = 199ns TO =200ns
.measure tran avgvall2bl244 AVG v(l2bl244) FROM = 199ns TO =200ns
.measure tran avgvall2bl245 AVG v(l2bl245) FROM = 199ns TO =200ns
.measure tran avgvall2bl246 AVG v(l2bl246) FROM = 199ns TO =200ns
.measure tran avgvall2bl247 AVG v(l2bl247) FROM = 199ns TO =200ns
.measure tran avgvall2bl248 AVG v(l2bl248) FROM = 199ns TO =200ns
.measure tran avgvall2bl249 AVG v(l2bl249) FROM = 199ns TO =200ns
.measure tran avgvall2bl250 AVG v(l2bl250) FROM = 199ns TO =200ns
.measure tran avgvall2bl251 AVG v(l2bl251) FROM = 199ns TO =200ns
.measure tran avgvall2bl252 AVG v(l2bl252) FROM = 199ns TO =200ns
.measure tran avgvall2bl253 AVG v(l2bl253) FROM = 199ns TO =200ns
.measure tran avgvall2bl254 AVG v(l2bl254) FROM = 199ns TO =200ns
.measure tran avgvall2bl255 AVG v(l2bl255) FROM = 199ns TO =200ns
.measure tran avgvall2bl256 AVG v(l2bl256) FROM = 199ns TO =200ns
.measure tran avgvall2bl257 AVG v(l2bl257) FROM = 199ns TO =200ns
.measure tran avgvall2bl258 AVG v(l2bl258) FROM = 199ns TO =200ns
.measure tran avgvall2bl259 AVG v(l2bl259) FROM = 199ns TO =200ns
.measure tran avgvall2bl260 AVG v(l2bl260) FROM = 199ns TO =200ns
.measure tran avgvall2bl261 AVG v(l2bl261) FROM = 199ns TO =200ns
.measure tran avgvall2bl262 AVG v(l2bl262) FROM = 199ns TO =200ns
.measure tran avgvall2bl263 AVG v(l2bl263) FROM = 199ns TO =200ns
.measure tran avgvall2bl264 AVG v(l2bl264) FROM = 199ns TO =200ns
.measure tran avgvall2bl265 AVG v(l2bl265) FROM = 199ns TO =200ns
.measure tran avgvall2bl266 AVG v(l2bl266) FROM = 199ns TO =200ns
.measure tran avgvall2bl267 AVG v(l2bl267) FROM = 199ns TO =200ns
.measure tran avgvall2bl268 AVG v(l2bl268) FROM = 199ns TO =200ns
.measure tran avgvall2bl269 AVG v(l2bl269) FROM = 199ns TO =200ns
.measure tran avgvall2bl270 AVG v(l2bl270) FROM = 199ns TO =200ns
.measure tran avgvall2bl271 AVG v(l2bl271) FROM = 199ns TO =200ns
.measure tran avgvall2bl272 AVG v(l2bl272) FROM = 199ns TO =200ns
.measure tran avgvall2bl273 AVG v(l2bl273) FROM = 199ns TO =200ns
.measure tran avgvall2bl274 AVG v(l2bl274) FROM = 199ns TO =200ns
.measure tran avgvall2bl275 AVG v(l2bl275) FROM = 199ns TO =200ns
.measure tran avgvall2bl276 AVG v(l2bl276) FROM = 199ns TO =200ns
.measure tran avgvall2bl277 AVG v(l2bl277) FROM = 199ns TO =200ns
.measure tran avgvall2bl278 AVG v(l2bl278) FROM = 199ns TO =200ns
.measure tran avgvall2bl279 AVG v(l2bl279) FROM = 199ns TO =200ns
.measure tran avgvall2bl280 AVG v(l2bl280) FROM = 199ns TO =200ns
.measure tran avgvall2bl281 AVG v(l2bl281) FROM = 199ns TO =200ns
.measure tran avgvall2bl282 AVG v(l2bl282) FROM = 199ns TO =200ns
.measure tran avgvall2bl283 AVG v(l2bl283) FROM = 199ns TO =200ns
.measure tran avgvall2bl284 AVG v(l2bl284) FROM = 199ns TO =200ns
.measure tran avgvall2bl285 AVG v(l2bl285) FROM = 199ns TO =200ns
.measure tran avgvall2bl286 AVG v(l2bl286) FROM = 199ns TO =200ns
.measure tran avgvall2bl287 AVG v(l2bl287) FROM = 199ns TO =200ns
.measure tran avgvall2bl288 AVG v(l2bl288) FROM = 199ns TO =200ns
.measure tran avgvall2bl289 AVG v(l2bl289) FROM = 199ns TO =200ns
.measure tran avgvall2bl290 AVG v(l2bl290) FROM = 199ns TO =200ns
.measure tran avgvall2bl291 AVG v(l2bl291) FROM = 199ns TO =200ns
.measure tran avgvall2bl292 AVG v(l2bl292) FROM = 199ns TO =200ns
.measure tran avgvall2bl293 AVG v(l2bl293) FROM = 199ns TO =200ns
.measure tran avgvall2bl294 AVG v(l2bl294) FROM = 199ns TO =200ns
.measure tran avgvall2bl295 AVG v(l2bl295) FROM = 199ns TO =200ns
.measure tran avgvall2bl296 AVG v(l2bl296) FROM = 199ns TO =200ns
.measure tran avgvall2bl297 AVG v(l2bl297) FROM = 199ns TO =200ns
.measure tran avgvall2bl298 AVG v(l2bl298) FROM = 199ns TO =200ns
.measure tran avgvall2bl299 AVG v(l2bl299) FROM = 199ns TO =200ns
.measure tran avgvall2bl300 AVG v(l2bl300) FROM = 199ns TO =200ns
.measure tran avgvall2bl301 AVG v(l2bl301) FROM = 199ns TO =200ns
.measure tran avgvall2bl302 AVG v(l2bl302) FROM = 199ns TO =200ns
.measure tran avgvall2bl303 AVG v(l2bl303) FROM = 199ns TO =200ns
.measure tran avgvall2bl304 AVG v(l2bl304) FROM = 199ns TO =200ns
.measure tran avgvall2bl305 AVG v(l2bl305) FROM = 199ns TO =200ns
.measure tran avgvall2bl306 AVG v(l2bl306) FROM = 199ns TO =200ns
.measure tran avgvall2bl307 AVG v(l2bl307) FROM = 199ns TO =200ns
.measure tran avgvall2bl308 AVG v(l2bl308) FROM = 199ns TO =200ns
.measure tran avgvall2bl309 AVG v(l2bl309) FROM = 199ns TO =200ns
.measure tran avgvall2bl310 AVG v(l2bl310) FROM = 199ns TO =200ns
.measure tran avgvall2bl311 AVG v(l2bl311) FROM = 199ns TO =200ns
.measure tran avgvall2bl312 AVG v(l2bl312) FROM = 199ns TO =200ns
.measure tran avgvall2bl313 AVG v(l2bl313) FROM = 199ns TO =200ns
.measure tran avgvall2bl314 AVG v(l2bl314) FROM = 199ns TO =200ns
.measure tran avgvall2bl315 AVG v(l2bl315) FROM = 199ns TO =200ns
.measure tran avgvall2bl316 AVG v(l2bl316) FROM = 199ns TO =200ns
.measure tran avgvall2bl317 AVG v(l2bl317) FROM = 199ns TO =200ns
.measure tran avgvall2bl318 AVG v(l2bl318) FROM = 199ns TO =200ns
.measure tran avgvall2bl319 AVG v(l2bl319) FROM = 199ns TO =200ns
.measure tran avgvall2bl320 AVG v(l2bl320) FROM = 199ns TO =200ns
.measure tran avgvall2bl321 AVG v(l2bl321) FROM = 199ns TO =200ns
.measure tran avgvall2bl322 AVG v(l2bl322) FROM = 199ns TO =200ns
.measure tran avgvall2bl323 AVG v(l2bl323) FROM = 199ns TO =200ns
.measure tran avgvall2bl324 AVG v(l2bl324) FROM = 199ns TO =200ns
.measure tran avgvall2bl325 AVG v(l2bl325) FROM = 199ns TO =200ns
.measure tran avgvall2bl326 AVG v(l2bl326) FROM = 199ns TO =200ns
.measure tran avgvall2bl327 AVG v(l2bl327) FROM = 199ns TO =200ns
.measure tran avgvall2bl328 AVG v(l2bl328) FROM = 199ns TO =200ns
.measure tran avgvall2bl329 AVG v(l2bl329) FROM = 199ns TO =200ns
.measure tran avgvall2bl330 AVG v(l2bl330) FROM = 199ns TO =200ns
.measure tran avgvall2bl331 AVG v(l2bl331) FROM = 199ns TO =200ns
.measure tran avgvall2bl332 AVG v(l2bl332) FROM = 199ns TO =200ns
.measure tran avgvall2bl333 AVG v(l2bl333) FROM = 199ns TO =200ns
.measure tran avgvall2bl334 AVG v(l2bl334) FROM = 199ns TO =200ns
.measure tran avgvall2bl335 AVG v(l2bl335) FROM = 199ns TO =200ns
.measure tran avgvall2bl336 AVG v(l2bl336) FROM = 199ns TO =200ns
.measure tran avgvall2bl337 AVG v(l2bl337) FROM = 199ns TO =200ns
.measure tran avgvall2bl338 AVG v(l2bl338) FROM = 199ns TO =200ns
.measure tran avgvall2bl339 AVG v(l2bl339) FROM = 199ns TO =200ns
.measure tran avgvall2bl340 AVG v(l2bl340) FROM = 199ns TO =200ns
.measure tran avgvall2bl341 AVG v(l2bl341) FROM = 199ns TO =200ns
.measure tran avgvall2bl342 AVG v(l2bl342) FROM = 199ns TO =200ns
.measure tran avgvall2bl343 AVG v(l2bl343) FROM = 199ns TO =200ns
.measure tran avgvall2bl344 AVG v(l2bl344) FROM = 199ns TO =200ns
.measure tran avgvall2bl345 AVG v(l2bl345) FROM = 199ns TO =200ns
.measure tran avgvall2bl346 AVG v(l2bl346) FROM = 199ns TO =200ns
.measure tran avgvall2bl347 AVG v(l2bl347) FROM = 199ns TO =200ns
.measure tran avgvall2bl348 AVG v(l2bl348) FROM = 199ns TO =200ns
.measure tran avgvall2bl349 AVG v(l2bl349) FROM = 199ns TO =200ns
.measure tran avgvall2bl350 AVG v(l2bl350) FROM = 199ns TO =200ns
.measure tran avgvall2bl351 AVG v(l2bl351) FROM = 199ns TO =200ns
.measure tran avgvall2bl352 AVG v(l2bl352) FROM = 199ns TO =200ns
.measure tran avgvall2bl353 AVG v(l2bl353) FROM = 199ns TO =200ns
.measure tran avgvall2bl354 AVG v(l2bl354) FROM = 199ns TO =200ns
.measure tran avgvall2bl355 AVG v(l2bl355) FROM = 199ns TO =200ns
.measure tran avgvall2bl356 AVG v(l2bl356) FROM = 199ns TO =200ns
.measure tran avgvall2bl357 AVG v(l2bl357) FROM = 199ns TO =200ns
.measure tran avgvall2bl358 AVG v(l2bl358) FROM = 199ns TO =200ns
.measure tran avgvall2bl359 AVG v(l2bl359) FROM = 199ns TO =200ns
.measure tran avgvall2bl360 AVG v(l2bl360) FROM = 199ns TO =200ns
.measure tran avgvall2bl361 AVG v(l2bl361) FROM = 199ns TO =200ns
.measure tran avgvall2bl362 AVG v(l2bl362) FROM = 199ns TO =200ns
.measure tran avgvall2bl363 AVG v(l2bl363) FROM = 199ns TO =200ns
.measure tran avgvall2bl364 AVG v(l2bl364) FROM = 199ns TO =200ns
.measure tran avgvall2bl365 AVG v(l2bl365) FROM = 199ns TO =200ns
.measure tran avgvall2bl366 AVG v(l2bl366) FROM = 199ns TO =200ns
.measure tran avgvall2bl367 AVG v(l2bl367) FROM = 199ns TO =200ns
.measure tran avgvall2bl368 AVG v(l2bl368) FROM = 199ns TO =200ns
.measure tran avgvall2bl369 AVG v(l2bl369) FROM = 199ns TO =200ns
.measure tran avgvall2bl370 AVG v(l2bl370) FROM = 199ns TO =200ns
.measure tran avgvall2bl371 AVG v(l2bl371) FROM = 199ns TO =200ns
.measure tran avgvall2bl372 AVG v(l2bl372) FROM = 199ns TO =200ns
.measure tran avgvall2bl373 AVG v(l2bl373) FROM = 199ns TO =200ns
.measure tran avgvall2bl374 AVG v(l2bl374) FROM = 199ns TO =200ns
.measure tran avgvall2bl375 AVG v(l2bl375) FROM = 199ns TO =200ns
.measure tran avgvall2bl376 AVG v(l2bl376) FROM = 199ns TO =200ns
.measure tran avgvall2bl377 AVG v(l2bl377) FROM = 199ns TO =200ns
.measure tran avgvall2bl378 AVG v(l2bl378) FROM = 199ns TO =200ns
.measure tran avgvall2bl379 AVG v(l2bl379) FROM = 199ns TO =200ns
.measure tran avgvall2bl380 AVG v(l2bl380) FROM = 199ns TO =200ns
.measure tran avgvall2bl381 AVG v(l2bl381) FROM = 199ns TO =200ns
.measure tran avgvall2bl382 AVG v(l2bl382) FROM = 199ns TO =200ns
.measure tran avgvall2bl383 AVG v(l2bl383) FROM = 199ns TO =200ns
.measure tran avgvall2bl384 AVG v(l2bl384) FROM = 199ns TO =200ns
.measure tran avgvall2bl385 AVG v(l2bl385) FROM = 199ns TO =200ns
.measure tran avgvall2bl386 AVG v(l2bl386) FROM = 199ns TO =200ns
.measure tran avgvall2bl387 AVG v(l2bl387) FROM = 199ns TO =200ns
.measure tran avgvall2bl388 AVG v(l2bl388) FROM = 199ns TO =200ns
.measure tran avgvall2bl389 AVG v(l2bl389) FROM = 199ns TO =200ns
.measure tran avgvall2bl390 AVG v(l2bl390) FROM = 199ns TO =200ns
.measure tran avgvall2bl391 AVG v(l2bl391) FROM = 199ns TO =200ns
.measure tran avgvall2bl392 AVG v(l2bl392) FROM = 199ns TO =200ns
.measure tran avgvall2bl393 AVG v(l2bl393) FROM = 199ns TO =200ns
.measure tran avgvall2bl394 AVG v(l2bl394) FROM = 199ns TO =200ns
.measure tran avgvall2bl395 AVG v(l2bl395) FROM = 199ns TO =200ns
.measure tran avgvall2bl396 AVG v(l2bl396) FROM = 199ns TO =200ns
.measure tran avgvall2bl397 AVG v(l2bl397) FROM = 199ns TO =200ns
.measure tran avgvall2bl398 AVG v(l2bl398) FROM = 199ns TO =200ns
.measure tran avgvall2bl399 AVG v(l2bl399) FROM = 199ns TO =200ns
.measure tran avgvall2bl400 AVG v(l2bl400) FROM = 199ns TO =200ns
.measure tran avgvall2bl401 AVG v(l2bl401) FROM = 199ns TO =200ns
.measure tran avgvall2bl402 AVG v(l2bl402) FROM = 199ns TO =200ns
.measure tran avgvall2bl403 AVG v(l2bl403) FROM = 199ns TO =200ns
.measure tran avgvall2bl404 AVG v(l2bl404) FROM = 199ns TO =200ns
.measure tran avgvall2bl405 AVG v(l2bl405) FROM = 199ns TO =200ns
.measure tran avgvall2bl406 AVG v(l2bl406) FROM = 199ns TO =200ns
.measure tran avgvall2bl407 AVG v(l2bl407) FROM = 199ns TO =200ns
.measure tran avgvall2bl408 AVG v(l2bl408) FROM = 199ns TO =200ns
.measure tran avgvall2bl409 AVG v(l2bl409) FROM = 199ns TO =200ns
.measure tran avgvall2bl410 AVG v(l2bl410) FROM = 199ns TO =200ns
.measure tran avgvall2bl411 AVG v(l2bl411) FROM = 199ns TO =200ns
.measure tran avgvall2bl412 AVG v(l2bl412) FROM = 199ns TO =200ns
.measure tran avgvall2bl413 AVG v(l2bl413) FROM = 199ns TO =200ns
.measure tran avgvall2bl414 AVG v(l2bl414) FROM = 199ns TO =200ns
.measure tran avgvall2bl415 AVG v(l2bl415) FROM = 199ns TO =200ns
.measure tran avgvall2bl416 AVG v(l2bl416) FROM = 199ns TO =200ns
.measure tran avgvall2bl417 AVG v(l2bl417) FROM = 199ns TO =200ns
.measure tran avgvall2bl418 AVG v(l2bl418) FROM = 199ns TO =200ns
.measure tran avgvall2bl419 AVG v(l2bl419) FROM = 199ns TO =200ns
.measure tran avgvall2bl420 AVG v(l2bl420) FROM = 199ns TO =200ns
.measure tran avgvall2bl421 AVG v(l2bl421) FROM = 199ns TO =200ns
.measure tran avgvall2bl422 AVG v(l2bl422) FROM = 199ns TO =200ns
.measure tran avgvall2bl423 AVG v(l2bl423) FROM = 199ns TO =200ns
.measure tran avgvall2bl424 AVG v(l2bl424) FROM = 199ns TO =200ns
.measure tran avgvall2bl425 AVG v(l2bl425) FROM = 199ns TO =200ns
.measure tran avgvall2bl426 AVG v(l2bl426) FROM = 199ns TO =200ns
.measure tran avgvall2bl427 AVG v(l2bl427) FROM = 199ns TO =200ns
.measure tran avgvall2bl428 AVG v(l2bl428) FROM = 199ns TO =200ns
.measure tran avgvall2bl429 AVG v(l2bl429) FROM = 199ns TO =200ns
.measure tran avgvall2bl430 AVG v(l2bl430) FROM = 199ns TO =200ns
.measure tran avgvall2bl431 AVG v(l2bl431) FROM = 199ns TO =200ns
.measure tran avgvall2bl432 AVG v(l2bl432) FROM = 199ns TO =200ns
.measure tran avgvall2bl433 AVG v(l2bl433) FROM = 199ns TO =200ns
.measure tran avgvall2bl434 AVG v(l2bl434) FROM = 199ns TO =200ns
.measure tran avgvall2bl435 AVG v(l2bl435) FROM = 199ns TO =200ns
.measure tran avgvall2bl436 AVG v(l2bl436) FROM = 199ns TO =200ns
.measure tran avgvall2bl437 AVG v(l2bl437) FROM = 199ns TO =200ns
.measure tran avgvall2bl438 AVG v(l2bl438) FROM = 199ns TO =200ns
.measure tran avgvall2bl439 AVG v(l2bl439) FROM = 199ns TO =200ns
.measure tran avgvall2bl440 AVG v(l2bl440) FROM = 199ns TO =200ns
.measure tran avgvall2bl441 AVG v(l2bl441) FROM = 199ns TO =200ns
.measure tran avgvall2bl442 AVG v(l2bl442) FROM = 199ns TO =200ns
.measure tran avgvall2bl443 AVG v(l2bl443) FROM = 199ns TO =200ns
.measure tran avgvall2bl444 AVG v(l2bl444) FROM = 199ns TO =200ns
.measure tran avgvall2bl445 AVG v(l2bl445) FROM = 199ns TO =200ns
.measure tran avgvall2bl446 AVG v(l2bl446) FROM = 199ns TO =200ns
.measure tran avgvall2bl447 AVG v(l2bl447) FROM = 199ns TO =200ns
.measure tran avgvall2bl448 AVG v(l2bl448) FROM = 199ns TO =200ns
.measure tran avgvall2bl449 AVG v(l2bl449) FROM = 199ns TO =200ns
.measure tran avgvall2bl450 AVG v(l2bl450) FROM = 199ns TO =200ns
.measure tran avgvall2bl451 AVG v(l2bl451) FROM = 199ns TO =200ns
.measure tran avgvall2bl452 AVG v(l2bl452) FROM = 199ns TO =200ns
.measure tran avgvall2bl453 AVG v(l2bl453) FROM = 199ns TO =200ns
.measure tran avgvall2bl454 AVG v(l2bl454) FROM = 199ns TO =200ns
.measure tran avgvall2bl455 AVG v(l2bl455) FROM = 199ns TO =200ns
.measure tran avgvall2bl456 AVG v(l2bl456) FROM = 199ns TO =200ns
.measure tran avgvall2bl457 AVG v(l2bl457) FROM = 199ns TO =200ns
.measure tran avgvall2bl458 AVG v(l2bl458) FROM = 199ns TO =200ns
.measure tran avgvall2bl459 AVG v(l2bl459) FROM = 199ns TO =200ns
.measure tran avgvall2bl460 AVG v(l2bl460) FROM = 199ns TO =200ns
.measure tran avgvall2bl461 AVG v(l2bl461) FROM = 199ns TO =200ns
.measure tran avgvall2bl462 AVG v(l2bl462) FROM = 199ns TO =200ns
.measure tran avgvall2bl463 AVG v(l2bl463) FROM = 199ns TO =200ns
.measure tran avgvall2bl464 AVG v(l2bl464) FROM = 199ns TO =200ns
.measure tran avgvall2bl465 AVG v(l2bl465) FROM = 199ns TO =200ns
.measure tran avgvall2bl466 AVG v(l2bl466) FROM = 199ns TO =200ns
.measure tran avgvall2bl467 AVG v(l2bl467) FROM = 199ns TO =200ns
.measure tran avgvall2bl468 AVG v(l2bl468) FROM = 199ns TO =200ns
.measure tran avgvall2bl469 AVG v(l2bl469) FROM = 199ns TO =200ns
.measure tran avgvall2bl470 AVG v(l2bl470) FROM = 199ns TO =200ns
.measure tran avgvall2bl471 AVG v(l2bl471) FROM = 199ns TO =200ns
.measure tran avgvall2bl472 AVG v(l2bl472) FROM = 199ns TO =200ns
.measure tran avgvall2bl473 AVG v(l2bl473) FROM = 199ns TO =200ns
.measure tran avgvall2bl474 AVG v(l2bl474) FROM = 199ns TO =200ns
.measure tran avgvall2bl475 AVG v(l2bl475) FROM = 199ns TO =200ns
.measure tran avgvall2bl476 AVG v(l2bl476) FROM = 199ns TO =200ns
.measure tran avgvall2bl477 AVG v(l2bl477) FROM = 199ns TO =200ns
.measure tran avgvall2bl478 AVG v(l2bl478) FROM = 199ns TO =200ns
.measure tran avgvall2bl479 AVG v(l2bl479) FROM = 199ns TO =200ns
.measure tran avgvall2bl480 AVG v(l2bl480) FROM = 199ns TO =200ns
.measure tran avgvall2bl481 AVG v(l2bl481) FROM = 199ns TO =200ns
.measure tran avgvall2bl482 AVG v(l2bl482) FROM = 199ns TO =200ns
.measure tran avgvall2bl483 AVG v(l2bl483) FROM = 199ns TO =200ns
.measure tran avgvall2bl484 AVG v(l2bl484) FROM = 199ns TO =200ns
.measure tran avgvall2bl485 AVG v(l2bl485) FROM = 199ns TO =200ns
.measure tran avgvall2bl486 AVG v(l2bl486) FROM = 199ns TO =200ns
.measure tran avgvall2bl487 AVG v(l2bl487) FROM = 199ns TO =200ns
.measure tran avgvall2bl488 AVG v(l2bl488) FROM = 199ns TO =200ns
.measure tran avgvall2bl489 AVG v(l2bl489) FROM = 199ns TO =200ns
.measure tran avgvall2bl490 AVG v(l2bl490) FROM = 199ns TO =200ns
.measure tran avgvall2bl491 AVG v(l2bl491) FROM = 199ns TO =200ns
.measure tran avgvall2bl492 AVG v(l2bl492) FROM = 199ns TO =200ns
.measure tran avgvall2bl493 AVG v(l2bl493) FROM = 199ns TO =200ns
.measure tran avgvall2bl494 AVG v(l2bl494) FROM = 199ns TO =200ns
.measure tran avgvall2bl495 AVG v(l2bl495) FROM = 199ns TO =200ns
.measure tran avgvall2bl496 AVG v(l2bl496) FROM = 199ns TO =200ns
.measure tran avgvall2bl497 AVG v(l2bl497) FROM = 199ns TO =200ns
.measure tran avgvall2bl498 AVG v(l2bl498) FROM = 199ns TO =200ns
.measure tran avgvall2bl499 AVG v(l2bl499) FROM = 199ns TO =200ns
.measure tran avgvall2bl500 AVG v(l2bl500) FROM = 199ns TO =200ns
.measure tran avgvall2bl501 AVG v(l2bl501) FROM = 199ns TO =200ns
.measure tran avgvall2bl502 AVG v(l2bl502) FROM = 199ns TO =200ns
.measure tran avgvall2bl503 AVG v(l2bl503) FROM = 199ns TO =200ns
.measure tran avgvall2bl504 AVG v(l2bl504) FROM = 199ns TO =200ns
.measure tran avgvall2bl505 AVG v(l2bl505) FROM = 199ns TO =200ns
.measure tran avgvall2bl506 AVG v(l2bl506) FROM = 199ns TO =200ns
.measure tran avgvall2bl507 AVG v(l2bl507) FROM = 199ns TO =200ns
.measure tran avgvall2bl508 AVG v(l2bl508) FROM = 199ns TO =200ns
.measure tran avgvall2bl509 AVG v(l2bl509) FROM = 199ns TO =200ns
.measure tran avgvall2bl510 AVG v(l2bl510) FROM = 199ns TO =200ns
.measure tran avgvall2bl511 AVG v(l2bl511) FROM = 199ns TO =200ns


.PROBE tran v(l3bl0)
.PROBE tran v(l3bl1)
.PROBE tran v(l3bl2)
.PROBE tran v(l3bl3)
.PROBE tran v(l3bl4)
.PROBE tran v(l3bl5)
.PROBE tran v(l3bl6)
.PROBE tran v(l3bl7)
.PROBE tran v(l3bl8)
.PROBE tran v(l3bl9)
.measure tran avgval0 AVG v(l3bl0) FROM = 199ns TO =200ns
.measure tran avgval1 AVG v(l3bl1) FROM = 199ns TO =200ns
.measure tran avgval2 AVG v(l3bl2) FROM = 199ns TO =200ns
.measure tran avgval3 AVG v(l3bl3) FROM = 199ns TO =200ns
.measure tran avgval4 AVG v(l3bl4) FROM = 199ns TO =200ns
.measure tran avgval5 AVG v(l3bl5) FROM = 199ns TO =200ns
.measure tran avgval6 AVG v(l3bl6) FROM = 199ns TO =200ns
.measure tran avgval7 AVG v(l3bl7) FROM = 199ns TO =200ns
.measure tran avgval8 AVG v(l3bl8) FROM = 199ns TO =200ns
.measure tran avgval9 AVG v(l3bl9) FROM = 199ns TO =200ns
.measure tran bld AVG v(bld) FROM = 99ns TO =100ns
.measure tran bldin AVG v(bldin) FROM = 99ns TO =100ns
.measure tran czabd AVG v(czabd) FROM = 99ns TO =100ns

.INCLUDE "/home/user68/design/rules/rohm180/spice/hspice/bu40n1.mdl"
.INCLUDE "/home/user68/DNN/insitu-training/20mv/bu40n3.mdl"
.LIB "/home/user68/design/rules/rohm180/spice/hspice/bu40n1.skw" NT
.LIB "/home/user68/design/rules/rohm180/spice/hspice/bu40n1.skw" PT

** Library name: reram
** Cell name: CELLD
** View name: schematic
.subckt CELLD bl sl wl wlb
m1 sl wlb net08 0 N L=180e-9 W=5e-6
m0 sl wl net09 0 N L=180e-9 W=5e-6
r1 net08 bl r1
r0 net09 bl r0
.ends CELLD
** End of subcircuit definition.

** Library name: reram
** Cell name: SAVM2
** View name: schematic
.subckt SAVM2 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N L=500e-9 W=3e-6
m2 net19 bl 0 0 N L=500e-9 W=3e-6
.ends SAVM2
** End of subcircuit definition.

** Library name: testRohm_n
** Cell name: INV1
** View name: schematic
.subckt INV1 g in out v
m1 out in v v P L=180e-9 W=5e-6
m0 out in g g N L=180e-9 W=2e-6
.ends INV1
** End of subcircuit definition.

** Library name: reram
** Cell name: CELLDREF
** View name: schematic
.subckt CELLDREF bl sl wl wlb
m1 sl wlb net13 net13 N L=180e-9 W=5e-6
m0 sl wl net14 net14 N L=180e-9 W=5e-6
r8 net018 bl 900e3
r7 net13 net018 10000e3
r6 net14 net020 900e3
r5 net020 bl 10000e3
r4 net017 bl 900e3
r3 net019 bl 10000e3
r1 net13 net017 10000e3
r0 net14 net019 900e3
.ends CELLDREF
** End of subcircuit definition.

** Library name: reram
** Cell name: XORNET4
** View name: schematic
.subckt SAVM2 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1602 L=500e-9 W=3e-6
m2 net19 bl 0 0 N2 L=500e-9 W=3e-6
.ends SAVM2

.subckt SAVM3 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1603 L=500e-9 W=3e-6
m2 net19 bl 0 0 N3 L=500e-9 W=3e-6
.ends SAVM3

.subckt SAVM4 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1604 L=500e-9 W=3e-6
m2 net19 bl 0 0 N4 L=500e-9 W=3e-6
.ends SAVM4

.subckt SAVM5 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1605 L=500e-9 W=3e-6
m2 net19 bl 0 0 N5 L=500e-9 W=3e-6
.ends SAVM5

.subckt SAVM6 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1606 L=500e-9 W=3e-6
m2 net19 bl 0 0 N6 L=500e-9 W=3e-6
.ends SAVM6

.subckt SAVM7 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1607 L=500e-9 W=3e-6
m2 net19 bl 0 0 N7 L=500e-9 W=3e-6
.ends SAVM7

.subckt SAVM8 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1608 L=500e-9 W=3e-6
m2 net19 bl 0 0 N8 L=500e-9 W=3e-6
.ends SAVM8

.subckt SAVM9 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1609 L=500e-9 W=3e-6
m2 net19 bl 0 0 N9 L=500e-9 W=3e-6
.ends SAVM9

.subckt SAVM10 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1610 L=500e-9 W=3e-6
m2 net19 bl 0 0 N10 L=500e-9 W=3e-6
.ends SAVM10

.subckt SAVM11 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1611 L=500e-9 W=3e-6
m2 net19 bl 0 0 N11 L=500e-9 W=3e-6
.ends SAVM11

.subckt SAVM12 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1612 L=500e-9 W=3e-6
m2 net19 bl 0 0 N12 L=500e-9 W=3e-6
.ends SAVM12

.subckt SAVM13 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1613 L=500e-9 W=3e-6
m2 net19 bl 0 0 N13 L=500e-9 W=3e-6
.ends SAVM13

.subckt SAVM14 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1614 L=500e-9 W=3e-6
m2 net19 bl 0 0 N14 L=500e-9 W=3e-6
.ends SAVM14

.subckt SAVM15 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1615 L=500e-9 W=3e-6
m2 net19 bl 0 0 N15 L=500e-9 W=3e-6
.ends SAVM15

.subckt SAVM16 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1616 L=500e-9 W=3e-6
m2 net19 bl 0 0 N16 L=500e-9 W=3e-6
.ends SAVM16

.subckt SAVM17 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1617 L=500e-9 W=3e-6
m2 net19 bl 0 0 N17 L=500e-9 W=3e-6
.ends SAVM17

.subckt SAVM18 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1618 L=500e-9 W=3e-6
m2 net19 bl 0 0 N18 L=500e-9 W=3e-6
.ends SAVM18

.subckt SAVM19 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1619 L=500e-9 W=3e-6
m2 net19 bl 0 0 N19 L=500e-9 W=3e-6
.ends SAVM19

.subckt SAVM20 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1620 L=500e-9 W=3e-6
m2 net19 bl 0 0 N20 L=500e-9 W=3e-6
.ends SAVM20

.subckt SAVM21 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1621 L=500e-9 W=3e-6
m2 net19 bl 0 0 N21 L=500e-9 W=3e-6
.ends SAVM21

.subckt SAVM22 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1622 L=500e-9 W=3e-6
m2 net19 bl 0 0 N22 L=500e-9 W=3e-6
.ends SAVM22

.subckt SAVM23 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1623 L=500e-9 W=3e-6
m2 net19 bl 0 0 N23 L=500e-9 W=3e-6
.ends SAVM23

.subckt SAVM24 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1624 L=500e-9 W=3e-6
m2 net19 bl 0 0 N24 L=500e-9 W=3e-6
.ends SAVM24

.subckt SAVM25 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1625 L=500e-9 W=3e-6
m2 net19 bl 0 0 N25 L=500e-9 W=3e-6
.ends SAVM25

.subckt SAVM26 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1626 L=500e-9 W=3e-6
m2 net19 bl 0 0 N26 L=500e-9 W=3e-6
.ends SAVM26

.subckt SAVM27 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1627 L=500e-9 W=3e-6
m2 net19 bl 0 0 N27 L=500e-9 W=3e-6
.ends SAVM27

.subckt SAVM28 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1628 L=500e-9 W=3e-6
m2 net19 bl 0 0 N28 L=500e-9 W=3e-6
.ends SAVM28

.subckt SAVM29 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1629 L=500e-9 W=3e-6
m2 net19 bl 0 0 N29 L=500e-9 W=3e-6
.ends SAVM29

.subckt SAVM30 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1630 L=500e-9 W=3e-6
m2 net19 bl 0 0 N30 L=500e-9 W=3e-6
.ends SAVM30

.subckt SAVM31 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1631 L=500e-9 W=3e-6
m2 net19 bl 0 0 N31 L=500e-9 W=3e-6
.ends SAVM31

.subckt SAVM32 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1632 L=500e-9 W=3e-6
m2 net19 bl 0 0 N32 L=500e-9 W=3e-6
.ends SAVM32

.subckt SAVM33 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1633 L=500e-9 W=3e-6
m2 net19 bl 0 0 N33 L=500e-9 W=3e-6
.ends SAVM33

.subckt SAVM34 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1634 L=500e-9 W=3e-6
m2 net19 bl 0 0 N34 L=500e-9 W=3e-6
.ends SAVM34

.subckt SAVM35 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1635 L=500e-9 W=3e-6
m2 net19 bl 0 0 N35 L=500e-9 W=3e-6
.ends SAVM35

.subckt SAVM36 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1636 L=500e-9 W=3e-6
m2 net19 bl 0 0 N36 L=500e-9 W=3e-6
.ends SAVM36

.subckt SAVM37 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1637 L=500e-9 W=3e-6
m2 net19 bl 0 0 N37 L=500e-9 W=3e-6
.ends SAVM37

.subckt SAVM38 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1638 L=500e-9 W=3e-6
m2 net19 bl 0 0 N38 L=500e-9 W=3e-6
.ends SAVM38

.subckt SAVM39 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1639 L=500e-9 W=3e-6
m2 net19 bl 0 0 N39 L=500e-9 W=3e-6
.ends SAVM39

.subckt SAVM40 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1640 L=500e-9 W=3e-6
m2 net19 bl 0 0 N40 L=500e-9 W=3e-6
.ends SAVM40

.subckt SAVM41 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1641 L=500e-9 W=3e-6
m2 net19 bl 0 0 N41 L=500e-9 W=3e-6
.ends SAVM41

.subckt SAVM42 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1642 L=500e-9 W=3e-6
m2 net19 bl 0 0 N42 L=500e-9 W=3e-6
.ends SAVM42

.subckt SAVM43 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1643 L=500e-9 W=3e-6
m2 net19 bl 0 0 N43 L=500e-9 W=3e-6
.ends SAVM43

.subckt SAVM44 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1644 L=500e-9 W=3e-6
m2 net19 bl 0 0 N44 L=500e-9 W=3e-6
.ends SAVM44

.subckt SAVM45 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1645 L=500e-9 W=3e-6
m2 net19 bl 0 0 N45 L=500e-9 W=3e-6
.ends SAVM45

.subckt SAVM46 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1646 L=500e-9 W=3e-6
m2 net19 bl 0 0 N46 L=500e-9 W=3e-6
.ends SAVM46

.subckt SAVM47 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1647 L=500e-9 W=3e-6
m2 net19 bl 0 0 N47 L=500e-9 W=3e-6
.ends SAVM47

.subckt SAVM48 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1648 L=500e-9 W=3e-6
m2 net19 bl 0 0 N48 L=500e-9 W=3e-6
.ends SAVM48

.subckt SAVM49 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1649 L=500e-9 W=3e-6
m2 net19 bl 0 0 N49 L=500e-9 W=3e-6
.ends SAVM49

.subckt SAVM50 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1650 L=500e-9 W=3e-6
m2 net19 bl 0 0 N50 L=500e-9 W=3e-6
.ends SAVM50

.subckt SAVM51 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1651 L=500e-9 W=3e-6
m2 net19 bl 0 0 N51 L=500e-9 W=3e-6
.ends SAVM51

.subckt SAVM52 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1652 L=500e-9 W=3e-6
m2 net19 bl 0 0 N52 L=500e-9 W=3e-6
.ends SAVM52

.subckt SAVM53 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1653 L=500e-9 W=3e-6
m2 net19 bl 0 0 N53 L=500e-9 W=3e-6
.ends SAVM53

.subckt SAVM54 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1654 L=500e-9 W=3e-6
m2 net19 bl 0 0 N54 L=500e-9 W=3e-6
.ends SAVM54

.subckt SAVM55 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1655 L=500e-9 W=3e-6
m2 net19 bl 0 0 N55 L=500e-9 W=3e-6
.ends SAVM55

.subckt SAVM56 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1656 L=500e-9 W=3e-6
m2 net19 bl 0 0 N56 L=500e-9 W=3e-6
.ends SAVM56

.subckt SAVM57 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1657 L=500e-9 W=3e-6
m2 net19 bl 0 0 N57 L=500e-9 W=3e-6
.ends SAVM57

.subckt SAVM58 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1658 L=500e-9 W=3e-6
m2 net19 bl 0 0 N58 L=500e-9 W=3e-6
.ends SAVM58

.subckt SAVM59 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1659 L=500e-9 W=3e-6
m2 net19 bl 0 0 N59 L=500e-9 W=3e-6
.ends SAVM59

.subckt SAVM60 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1660 L=500e-9 W=3e-6
m2 net19 bl 0 0 N60 L=500e-9 W=3e-6
.ends SAVM60

.subckt SAVM61 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1661 L=500e-9 W=3e-6
m2 net19 bl 0 0 N61 L=500e-9 W=3e-6
.ends SAVM61

.subckt SAVM62 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1662 L=500e-9 W=3e-6
m2 net19 bl 0 0 N62 L=500e-9 W=3e-6
.ends SAVM62

.subckt SAVM63 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1663 L=500e-9 W=3e-6
m2 net19 bl 0 0 N63 L=500e-9 W=3e-6
.ends SAVM63

.subckt SAVM64 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1664 L=500e-9 W=3e-6
m2 net19 bl 0 0 N64 L=500e-9 W=3e-6
.ends SAVM64

.subckt SAVM65 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1665 L=500e-9 W=3e-6
m2 net19 bl 0 0 N65 L=500e-9 W=3e-6
.ends SAVM65

.subckt SAVM66 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1666 L=500e-9 W=3e-6
m2 net19 bl 0 0 N66 L=500e-9 W=3e-6
.ends SAVM66

.subckt SAVM67 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1667 L=500e-9 W=3e-6
m2 net19 bl 0 0 N67 L=500e-9 W=3e-6
.ends SAVM67

.subckt SAVM68 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1668 L=500e-9 W=3e-6
m2 net19 bl 0 0 N68 L=500e-9 W=3e-6
.ends SAVM68

.subckt SAVM69 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1669 L=500e-9 W=3e-6
m2 net19 bl 0 0 N69 L=500e-9 W=3e-6
.ends SAVM69

.subckt SAVM70 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1670 L=500e-9 W=3e-6
m2 net19 bl 0 0 N70 L=500e-9 W=3e-6
.ends SAVM70

.subckt SAVM71 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1671 L=500e-9 W=3e-6
m2 net19 bl 0 0 N71 L=500e-9 W=3e-6
.ends SAVM71

.subckt SAVM72 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1672 L=500e-9 W=3e-6
m2 net19 bl 0 0 N72 L=500e-9 W=3e-6
.ends SAVM72

.subckt SAVM73 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1673 L=500e-9 W=3e-6
m2 net19 bl 0 0 N73 L=500e-9 W=3e-6
.ends SAVM73

.subckt SAVM74 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1674 L=500e-9 W=3e-6
m2 net19 bl 0 0 N74 L=500e-9 W=3e-6
.ends SAVM74

.subckt SAVM75 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1675 L=500e-9 W=3e-6
m2 net19 bl 0 0 N75 L=500e-9 W=3e-6
.ends SAVM75

.subckt SAVM76 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1676 L=500e-9 W=3e-6
m2 net19 bl 0 0 N76 L=500e-9 W=3e-6
.ends SAVM76

.subckt SAVM77 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1677 L=500e-9 W=3e-6
m2 net19 bl 0 0 N77 L=500e-9 W=3e-6
.ends SAVM77

.subckt SAVM78 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1678 L=500e-9 W=3e-6
m2 net19 bl 0 0 N78 L=500e-9 W=3e-6
.ends SAVM78

.subckt SAVM79 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1679 L=500e-9 W=3e-6
m2 net19 bl 0 0 N79 L=500e-9 W=3e-6
.ends SAVM79

.subckt SAVM80 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1680 L=500e-9 W=3e-6
m2 net19 bl 0 0 N80 L=500e-9 W=3e-6
.ends SAVM80

.subckt SAVM81 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1681 L=500e-9 W=3e-6
m2 net19 bl 0 0 N81 L=500e-9 W=3e-6
.ends SAVM81

.subckt SAVM82 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1682 L=500e-9 W=3e-6
m2 net19 bl 0 0 N82 L=500e-9 W=3e-6
.ends SAVM82

.subckt SAVM83 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1683 L=500e-9 W=3e-6
m2 net19 bl 0 0 N83 L=500e-9 W=3e-6
.ends SAVM83

.subckt SAVM84 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1684 L=500e-9 W=3e-6
m2 net19 bl 0 0 N84 L=500e-9 W=3e-6
.ends SAVM84

.subckt SAVM85 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1685 L=500e-9 W=3e-6
m2 net19 bl 0 0 N85 L=500e-9 W=3e-6
.ends SAVM85

.subckt SAVM86 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1686 L=500e-9 W=3e-6
m2 net19 bl 0 0 N86 L=500e-9 W=3e-6
.ends SAVM86

.subckt SAVM87 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1687 L=500e-9 W=3e-6
m2 net19 bl 0 0 N87 L=500e-9 W=3e-6
.ends SAVM87

.subckt SAVM88 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1688 L=500e-9 W=3e-6
m2 net19 bl 0 0 N88 L=500e-9 W=3e-6
.ends SAVM88

.subckt SAVM89 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1689 L=500e-9 W=3e-6
m2 net19 bl 0 0 N89 L=500e-9 W=3e-6
.ends SAVM89

.subckt SAVM90 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1690 L=500e-9 W=3e-6
m2 net19 bl 0 0 N90 L=500e-9 W=3e-6
.ends SAVM90

.subckt SAVM91 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1691 L=500e-9 W=3e-6
m2 net19 bl 0 0 N91 L=500e-9 W=3e-6
.ends SAVM91

.subckt SAVM92 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1692 L=500e-9 W=3e-6
m2 net19 bl 0 0 N92 L=500e-9 W=3e-6
.ends SAVM92

.subckt SAVM93 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1693 L=500e-9 W=3e-6
m2 net19 bl 0 0 N93 L=500e-9 W=3e-6
.ends SAVM93

.subckt SAVM94 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1694 L=500e-9 W=3e-6
m2 net19 bl 0 0 N94 L=500e-9 W=3e-6
.ends SAVM94

.subckt SAVM95 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1695 L=500e-9 W=3e-6
m2 net19 bl 0 0 N95 L=500e-9 W=3e-6
.ends SAVM95

.subckt SAVM96 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1696 L=500e-9 W=3e-6
m2 net19 bl 0 0 N96 L=500e-9 W=3e-6
.ends SAVM96

.subckt SAVM97 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1697 L=500e-9 W=3e-6
m2 net19 bl 0 0 N97 L=500e-9 W=3e-6
.ends SAVM97

.subckt SAVM98 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1698 L=500e-9 W=3e-6
m2 net19 bl 0 0 N98 L=500e-9 W=3e-6
.ends SAVM98

.subckt SAVM99 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1699 L=500e-9 W=3e-6
m2 net19 bl 0 0 N99 L=500e-9 W=3e-6
.ends SAVM99

.subckt SAVM100 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1700 L=500e-9 W=3e-6
m2 net19 bl 0 0 N100 L=500e-9 W=3e-6
.ends SAVM100

.subckt SAVM101 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1701 L=500e-9 W=3e-6
m2 net19 bl 0 0 N101 L=500e-9 W=3e-6
.ends SAVM101

.subckt SAVM102 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1702 L=500e-9 W=3e-6
m2 net19 bl 0 0 N102 L=500e-9 W=3e-6
.ends SAVM102

.subckt SAVM103 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1703 L=500e-9 W=3e-6
m2 net19 bl 0 0 N103 L=500e-9 W=3e-6
.ends SAVM103

.subckt SAVM104 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1704 L=500e-9 W=3e-6
m2 net19 bl 0 0 N104 L=500e-9 W=3e-6
.ends SAVM104

.subckt SAVM105 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1705 L=500e-9 W=3e-6
m2 net19 bl 0 0 N105 L=500e-9 W=3e-6
.ends SAVM105

.subckt SAVM106 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1706 L=500e-9 W=3e-6
m2 net19 bl 0 0 N106 L=500e-9 W=3e-6
.ends SAVM106

.subckt SAVM107 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1707 L=500e-9 W=3e-6
m2 net19 bl 0 0 N107 L=500e-9 W=3e-6
.ends SAVM107

.subckt SAVM108 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1708 L=500e-9 W=3e-6
m2 net19 bl 0 0 N108 L=500e-9 W=3e-6
.ends SAVM108

.subckt SAVM109 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1709 L=500e-9 W=3e-6
m2 net19 bl 0 0 N109 L=500e-9 W=3e-6
.ends SAVM109

.subckt SAVM110 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1710 L=500e-9 W=3e-6
m2 net19 bl 0 0 N110 L=500e-9 W=3e-6
.ends SAVM110

.subckt SAVM111 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1711 L=500e-9 W=3e-6
m2 net19 bl 0 0 N111 L=500e-9 W=3e-6
.ends SAVM111

.subckt SAVM112 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1712 L=500e-9 W=3e-6
m2 net19 bl 0 0 N112 L=500e-9 W=3e-6
.ends SAVM112

.subckt SAVM113 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1713 L=500e-9 W=3e-6
m2 net19 bl 0 0 N113 L=500e-9 W=3e-6
.ends SAVM113

.subckt SAVM114 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1714 L=500e-9 W=3e-6
m2 net19 bl 0 0 N114 L=500e-9 W=3e-6
.ends SAVM114

.subckt SAVM115 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1715 L=500e-9 W=3e-6
m2 net19 bl 0 0 N115 L=500e-9 W=3e-6
.ends SAVM115

.subckt SAVM116 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1716 L=500e-9 W=3e-6
m2 net19 bl 0 0 N116 L=500e-9 W=3e-6
.ends SAVM116

.subckt SAVM117 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1717 L=500e-9 W=3e-6
m2 net19 bl 0 0 N117 L=500e-9 W=3e-6
.ends SAVM117

.subckt SAVM118 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1718 L=500e-9 W=3e-6
m2 net19 bl 0 0 N118 L=500e-9 W=3e-6
.ends SAVM118

.subckt SAVM119 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1719 L=500e-9 W=3e-6
m2 net19 bl 0 0 N119 L=500e-9 W=3e-6
.ends SAVM119

.subckt SAVM120 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1720 L=500e-9 W=3e-6
m2 net19 bl 0 0 N120 L=500e-9 W=3e-6
.ends SAVM120

.subckt SAVM121 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1721 L=500e-9 W=3e-6
m2 net19 bl 0 0 N121 L=500e-9 W=3e-6
.ends SAVM121

.subckt SAVM122 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1722 L=500e-9 W=3e-6
m2 net19 bl 0 0 N122 L=500e-9 W=3e-6
.ends SAVM122

.subckt SAVM123 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1723 L=500e-9 W=3e-6
m2 net19 bl 0 0 N123 L=500e-9 W=3e-6
.ends SAVM123

.subckt SAVM124 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1724 L=500e-9 W=3e-6
m2 net19 bl 0 0 N124 L=500e-9 W=3e-6
.ends SAVM124

.subckt SAVM125 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1725 L=500e-9 W=3e-6
m2 net19 bl 0 0 N125 L=500e-9 W=3e-6
.ends SAVM125

.subckt SAVM126 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1726 L=500e-9 W=3e-6
m2 net19 bl 0 0 N126 L=500e-9 W=3e-6
.ends SAVM126

.subckt SAVM127 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1727 L=500e-9 W=3e-6
m2 net19 bl 0 0 N127 L=500e-9 W=3e-6
.ends SAVM127

.subckt SAVM128 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1728 L=500e-9 W=3e-6
m2 net19 bl 0 0 N128 L=500e-9 W=3e-6
.ends SAVM128

.subckt SAVM129 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1729 L=500e-9 W=3e-6
m2 net19 bl 0 0 N129 L=500e-9 W=3e-6
.ends SAVM129

.subckt SAVM130 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1730 L=500e-9 W=3e-6
m2 net19 bl 0 0 N130 L=500e-9 W=3e-6
.ends SAVM130

.subckt SAVM131 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1731 L=500e-9 W=3e-6
m2 net19 bl 0 0 N131 L=500e-9 W=3e-6
.ends SAVM131

.subckt SAVM132 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1732 L=500e-9 W=3e-6
m2 net19 bl 0 0 N132 L=500e-9 W=3e-6
.ends SAVM132

.subckt SAVM133 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1733 L=500e-9 W=3e-6
m2 net19 bl 0 0 N133 L=500e-9 W=3e-6
.ends SAVM133

.subckt SAVM134 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1734 L=500e-9 W=3e-6
m2 net19 bl 0 0 N134 L=500e-9 W=3e-6
.ends SAVM134

.subckt SAVM135 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1735 L=500e-9 W=3e-6
m2 net19 bl 0 0 N135 L=500e-9 W=3e-6
.ends SAVM135

.subckt SAVM136 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1736 L=500e-9 W=3e-6
m2 net19 bl 0 0 N136 L=500e-9 W=3e-6
.ends SAVM136

.subckt SAVM137 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1737 L=500e-9 W=3e-6
m2 net19 bl 0 0 N137 L=500e-9 W=3e-6
.ends SAVM137

.subckt SAVM138 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1738 L=500e-9 W=3e-6
m2 net19 bl 0 0 N138 L=500e-9 W=3e-6
.ends SAVM138

.subckt SAVM139 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1739 L=500e-9 W=3e-6
m2 net19 bl 0 0 N139 L=500e-9 W=3e-6
.ends SAVM139

.subckt SAVM140 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1740 L=500e-9 W=3e-6
m2 net19 bl 0 0 N140 L=500e-9 W=3e-6
.ends SAVM140

.subckt SAVM141 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1741 L=500e-9 W=3e-6
m2 net19 bl 0 0 N141 L=500e-9 W=3e-6
.ends SAVM141

.subckt SAVM142 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1742 L=500e-9 W=3e-6
m2 net19 bl 0 0 N142 L=500e-9 W=3e-6
.ends SAVM142

.subckt SAVM143 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1743 L=500e-9 W=3e-6
m2 net19 bl 0 0 N143 L=500e-9 W=3e-6
.ends SAVM143

.subckt SAVM144 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1744 L=500e-9 W=3e-6
m2 net19 bl 0 0 N144 L=500e-9 W=3e-6
.ends SAVM144

.subckt SAVM145 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1745 L=500e-9 W=3e-6
m2 net19 bl 0 0 N145 L=500e-9 W=3e-6
.ends SAVM145

.subckt SAVM146 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1746 L=500e-9 W=3e-6
m2 net19 bl 0 0 N146 L=500e-9 W=3e-6
.ends SAVM146

.subckt SAVM147 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1747 L=500e-9 W=3e-6
m2 net19 bl 0 0 N147 L=500e-9 W=3e-6
.ends SAVM147

.subckt SAVM148 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1748 L=500e-9 W=3e-6
m2 net19 bl 0 0 N148 L=500e-9 W=3e-6
.ends SAVM148

.subckt SAVM149 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1749 L=500e-9 W=3e-6
m2 net19 bl 0 0 N149 L=500e-9 W=3e-6
.ends SAVM149

.subckt SAVM150 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1750 L=500e-9 W=3e-6
m2 net19 bl 0 0 N150 L=500e-9 W=3e-6
.ends SAVM150

.subckt SAVM151 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1751 L=500e-9 W=3e-6
m2 net19 bl 0 0 N151 L=500e-9 W=3e-6
.ends SAVM151

.subckt SAVM152 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1752 L=500e-9 W=3e-6
m2 net19 bl 0 0 N152 L=500e-9 W=3e-6
.ends SAVM152

.subckt SAVM153 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1753 L=500e-9 W=3e-6
m2 net19 bl 0 0 N153 L=500e-9 W=3e-6
.ends SAVM153

.subckt SAVM154 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1754 L=500e-9 W=3e-6
m2 net19 bl 0 0 N154 L=500e-9 W=3e-6
.ends SAVM154

.subckt SAVM155 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1755 L=500e-9 W=3e-6
m2 net19 bl 0 0 N155 L=500e-9 W=3e-6
.ends SAVM155

.subckt SAVM156 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1756 L=500e-9 W=3e-6
m2 net19 bl 0 0 N156 L=500e-9 W=3e-6
.ends SAVM156

.subckt SAVM157 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1757 L=500e-9 W=3e-6
m2 net19 bl 0 0 N157 L=500e-9 W=3e-6
.ends SAVM157

.subckt SAVM158 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1758 L=500e-9 W=3e-6
m2 net19 bl 0 0 N158 L=500e-9 W=3e-6
.ends SAVM158

.subckt SAVM159 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1759 L=500e-9 W=3e-6
m2 net19 bl 0 0 N159 L=500e-9 W=3e-6
.ends SAVM159

.subckt SAVM160 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1760 L=500e-9 W=3e-6
m2 net19 bl 0 0 N160 L=500e-9 W=3e-6
.ends SAVM160

.subckt SAVM161 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1761 L=500e-9 W=3e-6
m2 net19 bl 0 0 N161 L=500e-9 W=3e-6
.ends SAVM161

.subckt SAVM162 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1762 L=500e-9 W=3e-6
m2 net19 bl 0 0 N162 L=500e-9 W=3e-6
.ends SAVM162

.subckt SAVM163 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1763 L=500e-9 W=3e-6
m2 net19 bl 0 0 N163 L=500e-9 W=3e-6
.ends SAVM163

.subckt SAVM164 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1764 L=500e-9 W=3e-6
m2 net19 bl 0 0 N164 L=500e-9 W=3e-6
.ends SAVM164

.subckt SAVM165 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1765 L=500e-9 W=3e-6
m2 net19 bl 0 0 N165 L=500e-9 W=3e-6
.ends SAVM165

.subckt SAVM166 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1766 L=500e-9 W=3e-6
m2 net19 bl 0 0 N166 L=500e-9 W=3e-6
.ends SAVM166

.subckt SAVM167 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1767 L=500e-9 W=3e-6
m2 net19 bl 0 0 N167 L=500e-9 W=3e-6
.ends SAVM167

.subckt SAVM168 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1768 L=500e-9 W=3e-6
m2 net19 bl 0 0 N168 L=500e-9 W=3e-6
.ends SAVM168

.subckt SAVM169 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1769 L=500e-9 W=3e-6
m2 net19 bl 0 0 N169 L=500e-9 W=3e-6
.ends SAVM169

.subckt SAVM170 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1770 L=500e-9 W=3e-6
m2 net19 bl 0 0 N170 L=500e-9 W=3e-6
.ends SAVM170

.subckt SAVM171 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1771 L=500e-9 W=3e-6
m2 net19 bl 0 0 N171 L=500e-9 W=3e-6
.ends SAVM171

.subckt SAVM172 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1772 L=500e-9 W=3e-6
m2 net19 bl 0 0 N172 L=500e-9 W=3e-6
.ends SAVM172

.subckt SAVM173 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1773 L=500e-9 W=3e-6
m2 net19 bl 0 0 N173 L=500e-9 W=3e-6
.ends SAVM173

.subckt SAVM174 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1774 L=500e-9 W=3e-6
m2 net19 bl 0 0 N174 L=500e-9 W=3e-6
.ends SAVM174

.subckt SAVM175 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1775 L=500e-9 W=3e-6
m2 net19 bl 0 0 N175 L=500e-9 W=3e-6
.ends SAVM175

.subckt SAVM176 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1776 L=500e-9 W=3e-6
m2 net19 bl 0 0 N176 L=500e-9 W=3e-6
.ends SAVM176

.subckt SAVM177 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1777 L=500e-9 W=3e-6
m2 net19 bl 0 0 N177 L=500e-9 W=3e-6
.ends SAVM177

.subckt SAVM178 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1778 L=500e-9 W=3e-6
m2 net19 bl 0 0 N178 L=500e-9 W=3e-6
.ends SAVM178

.subckt SAVM179 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1779 L=500e-9 W=3e-6
m2 net19 bl 0 0 N179 L=500e-9 W=3e-6
.ends SAVM179

.subckt SAVM180 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1780 L=500e-9 W=3e-6
m2 net19 bl 0 0 N180 L=500e-9 W=3e-6
.ends SAVM180

.subckt SAVM181 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1781 L=500e-9 W=3e-6
m2 net19 bl 0 0 N181 L=500e-9 W=3e-6
.ends SAVM181

.subckt SAVM182 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1782 L=500e-9 W=3e-6
m2 net19 bl 0 0 N182 L=500e-9 W=3e-6
.ends SAVM182

.subckt SAVM183 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1783 L=500e-9 W=3e-6
m2 net19 bl 0 0 N183 L=500e-9 W=3e-6
.ends SAVM183

.subckt SAVM184 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1784 L=500e-9 W=3e-6
m2 net19 bl 0 0 N184 L=500e-9 W=3e-6
.ends SAVM184

.subckt SAVM185 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1785 L=500e-9 W=3e-6
m2 net19 bl 0 0 N185 L=500e-9 W=3e-6
.ends SAVM185

.subckt SAVM186 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1786 L=500e-9 W=3e-6
m2 net19 bl 0 0 N186 L=500e-9 W=3e-6
.ends SAVM186

.subckt SAVM187 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1787 L=500e-9 W=3e-6
m2 net19 bl 0 0 N187 L=500e-9 W=3e-6
.ends SAVM187

.subckt SAVM188 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1788 L=500e-9 W=3e-6
m2 net19 bl 0 0 N188 L=500e-9 W=3e-6
.ends SAVM188

.subckt SAVM189 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1789 L=500e-9 W=3e-6
m2 net19 bl 0 0 N189 L=500e-9 W=3e-6
.ends SAVM189

.subckt SAVM190 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1790 L=500e-9 W=3e-6
m2 net19 bl 0 0 N190 L=500e-9 W=3e-6
.ends SAVM190

.subckt SAVM191 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1791 L=500e-9 W=3e-6
m2 net19 bl 0 0 N191 L=500e-9 W=3e-6
.ends SAVM191

.subckt SAVM192 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1792 L=500e-9 W=3e-6
m2 net19 bl 0 0 N192 L=500e-9 W=3e-6
.ends SAVM192

.subckt SAVM193 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1793 L=500e-9 W=3e-6
m2 net19 bl 0 0 N193 L=500e-9 W=3e-6
.ends SAVM193

.subckt SAVM194 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1794 L=500e-9 W=3e-6
m2 net19 bl 0 0 N194 L=500e-9 W=3e-6
.ends SAVM194

.subckt SAVM195 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1795 L=500e-9 W=3e-6
m2 net19 bl 0 0 N195 L=500e-9 W=3e-6
.ends SAVM195

.subckt SAVM196 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1796 L=500e-9 W=3e-6
m2 net19 bl 0 0 N196 L=500e-9 W=3e-6
.ends SAVM196

.subckt SAVM197 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1797 L=500e-9 W=3e-6
m2 net19 bl 0 0 N197 L=500e-9 W=3e-6
.ends SAVM197

.subckt SAVM198 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1798 L=500e-9 W=3e-6
m2 net19 bl 0 0 N198 L=500e-9 W=3e-6
.ends SAVM198

.subckt SAVM199 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1799 L=500e-9 W=3e-6
m2 net19 bl 0 0 N199 L=500e-9 W=3e-6
.ends SAVM199

.subckt SAVM200 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1800 L=500e-9 W=3e-6
m2 net19 bl 0 0 N200 L=500e-9 W=3e-6
.ends SAVM200

.subckt SAVM201 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1801 L=500e-9 W=3e-6
m2 net19 bl 0 0 N201 L=500e-9 W=3e-6
.ends SAVM201

.subckt SAVM202 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1802 L=500e-9 W=3e-6
m2 net19 bl 0 0 N202 L=500e-9 W=3e-6
.ends SAVM202

.subckt SAVM203 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1803 L=500e-9 W=3e-6
m2 net19 bl 0 0 N203 L=500e-9 W=3e-6
.ends SAVM203

.subckt SAVM204 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1804 L=500e-9 W=3e-6
m2 net19 bl 0 0 N204 L=500e-9 W=3e-6
.ends SAVM204

.subckt SAVM205 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1805 L=500e-9 W=3e-6
m2 net19 bl 0 0 N205 L=500e-9 W=3e-6
.ends SAVM205

.subckt SAVM206 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1806 L=500e-9 W=3e-6
m2 net19 bl 0 0 N206 L=500e-9 W=3e-6
.ends SAVM206

.subckt SAVM207 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1807 L=500e-9 W=3e-6
m2 net19 bl 0 0 N207 L=500e-9 W=3e-6
.ends SAVM207

.subckt SAVM208 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1808 L=500e-9 W=3e-6
m2 net19 bl 0 0 N208 L=500e-9 W=3e-6
.ends SAVM208

.subckt SAVM209 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1809 L=500e-9 W=3e-6
m2 net19 bl 0 0 N209 L=500e-9 W=3e-6
.ends SAVM209

.subckt SAVM210 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1810 L=500e-9 W=3e-6
m2 net19 bl 0 0 N210 L=500e-9 W=3e-6
.ends SAVM210

.subckt SAVM211 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1811 L=500e-9 W=3e-6
m2 net19 bl 0 0 N211 L=500e-9 W=3e-6
.ends SAVM211

.subckt SAVM212 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1812 L=500e-9 W=3e-6
m2 net19 bl 0 0 N212 L=500e-9 W=3e-6
.ends SAVM212

.subckt SAVM213 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1813 L=500e-9 W=3e-6
m2 net19 bl 0 0 N213 L=500e-9 W=3e-6
.ends SAVM213

.subckt SAVM214 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1814 L=500e-9 W=3e-6
m2 net19 bl 0 0 N214 L=500e-9 W=3e-6
.ends SAVM214

.subckt SAVM215 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1815 L=500e-9 W=3e-6
m2 net19 bl 0 0 N215 L=500e-9 W=3e-6
.ends SAVM215

.subckt SAVM216 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1816 L=500e-9 W=3e-6
m2 net19 bl 0 0 N216 L=500e-9 W=3e-6
.ends SAVM216

.subckt SAVM217 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1817 L=500e-9 W=3e-6
m2 net19 bl 0 0 N217 L=500e-9 W=3e-6
.ends SAVM217

.subckt SAVM218 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1818 L=500e-9 W=3e-6
m2 net19 bl 0 0 N218 L=500e-9 W=3e-6
.ends SAVM218

.subckt SAVM219 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1819 L=500e-9 W=3e-6
m2 net19 bl 0 0 N219 L=500e-9 W=3e-6
.ends SAVM219

.subckt SAVM220 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1820 L=500e-9 W=3e-6
m2 net19 bl 0 0 N220 L=500e-9 W=3e-6
.ends SAVM220

.subckt SAVM221 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1821 L=500e-9 W=3e-6
m2 net19 bl 0 0 N221 L=500e-9 W=3e-6
.ends SAVM221

.subckt SAVM222 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1822 L=500e-9 W=3e-6
m2 net19 bl 0 0 N222 L=500e-9 W=3e-6
.ends SAVM222

.subckt SAVM223 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1823 L=500e-9 W=3e-6
m2 net19 bl 0 0 N223 L=500e-9 W=3e-6
.ends SAVM223

.subckt SAVM224 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1824 L=500e-9 W=3e-6
m2 net19 bl 0 0 N224 L=500e-9 W=3e-6
.ends SAVM224

.subckt SAVM225 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1825 L=500e-9 W=3e-6
m2 net19 bl 0 0 N225 L=500e-9 W=3e-6
.ends SAVM225

.subckt SAVM226 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1826 L=500e-9 W=3e-6
m2 net19 bl 0 0 N226 L=500e-9 W=3e-6
.ends SAVM226

.subckt SAVM227 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1827 L=500e-9 W=3e-6
m2 net19 bl 0 0 N227 L=500e-9 W=3e-6
.ends SAVM227

.subckt SAVM228 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1828 L=500e-9 W=3e-6
m2 net19 bl 0 0 N228 L=500e-9 W=3e-6
.ends SAVM228

.subckt SAVM229 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1829 L=500e-9 W=3e-6
m2 net19 bl 0 0 N229 L=500e-9 W=3e-6
.ends SAVM229

.subckt SAVM230 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1830 L=500e-9 W=3e-6
m2 net19 bl 0 0 N230 L=500e-9 W=3e-6
.ends SAVM230

.subckt SAVM231 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1831 L=500e-9 W=3e-6
m2 net19 bl 0 0 N231 L=500e-9 W=3e-6
.ends SAVM231

.subckt SAVM232 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1832 L=500e-9 W=3e-6
m2 net19 bl 0 0 N232 L=500e-9 W=3e-6
.ends SAVM232

.subckt SAVM233 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1833 L=500e-9 W=3e-6
m2 net19 bl 0 0 N233 L=500e-9 W=3e-6
.ends SAVM233

.subckt SAVM234 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1834 L=500e-9 W=3e-6
m2 net19 bl 0 0 N234 L=500e-9 W=3e-6
.ends SAVM234

.subckt SAVM235 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1835 L=500e-9 W=3e-6
m2 net19 bl 0 0 N235 L=500e-9 W=3e-6
.ends SAVM235

.subckt SAVM236 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1836 L=500e-9 W=3e-6
m2 net19 bl 0 0 N236 L=500e-9 W=3e-6
.ends SAVM236

.subckt SAVM237 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1837 L=500e-9 W=3e-6
m2 net19 bl 0 0 N237 L=500e-9 W=3e-6
.ends SAVM237

.subckt SAVM238 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1838 L=500e-9 W=3e-6
m2 net19 bl 0 0 N238 L=500e-9 W=3e-6
.ends SAVM238

.subckt SAVM239 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1839 L=500e-9 W=3e-6
m2 net19 bl 0 0 N239 L=500e-9 W=3e-6
.ends SAVM239

.subckt SAVM240 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1840 L=500e-9 W=3e-6
m2 net19 bl 0 0 N240 L=500e-9 W=3e-6
.ends SAVM240

.subckt SAVM241 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1841 L=500e-9 W=3e-6
m2 net19 bl 0 0 N241 L=500e-9 W=3e-6
.ends SAVM241

.subckt SAVM242 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1842 L=500e-9 W=3e-6
m2 net19 bl 0 0 N242 L=500e-9 W=3e-6
.ends SAVM242

.subckt SAVM243 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1843 L=500e-9 W=3e-6
m2 net19 bl 0 0 N243 L=500e-9 W=3e-6
.ends SAVM243

.subckt SAVM244 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1844 L=500e-9 W=3e-6
m2 net19 bl 0 0 N244 L=500e-9 W=3e-6
.ends SAVM244

.subckt SAVM245 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1845 L=500e-9 W=3e-6
m2 net19 bl 0 0 N245 L=500e-9 W=3e-6
.ends SAVM245

.subckt SAVM246 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1846 L=500e-9 W=3e-6
m2 net19 bl 0 0 N246 L=500e-9 W=3e-6
.ends SAVM246

.subckt SAVM247 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1847 L=500e-9 W=3e-6
m2 net19 bl 0 0 N247 L=500e-9 W=3e-6
.ends SAVM247

.subckt SAVM248 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1848 L=500e-9 W=3e-6
m2 net19 bl 0 0 N248 L=500e-9 W=3e-6
.ends SAVM248

.subckt SAVM249 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1849 L=500e-9 W=3e-6
m2 net19 bl 0 0 N249 L=500e-9 W=3e-6
.ends SAVM249

.subckt SAVM250 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1850 L=500e-9 W=3e-6
m2 net19 bl 0 0 N250 L=500e-9 W=3e-6
.ends SAVM250

.subckt SAVM251 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1851 L=500e-9 W=3e-6
m2 net19 bl 0 0 N251 L=500e-9 W=3e-6
.ends SAVM251

.subckt SAVM252 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1852 L=500e-9 W=3e-6
m2 net19 bl 0 0 N252 L=500e-9 W=3e-6
.ends SAVM252

.subckt SAVM253 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1853 L=500e-9 W=3e-6
m2 net19 bl 0 0 N253 L=500e-9 W=3e-6
.ends SAVM253

.subckt SAVM254 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1854 L=500e-9 W=3e-6
m2 net19 bl 0 0 N254 L=500e-9 W=3e-6
.ends SAVM254

.subckt SAVM255 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1855 L=500e-9 W=3e-6
m2 net19 bl 0 0 N255 L=500e-9 W=3e-6
.ends SAVM255

.subckt SAVM256 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1856 L=500e-9 W=3e-6
m2 net19 bl 0 0 N256 L=500e-9 W=3e-6
.ends SAVM256

.subckt SAVM257 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1857 L=500e-9 W=3e-6
m2 net19 bl 0 0 N257 L=500e-9 W=3e-6
.ends SAVM257

.subckt SAVM258 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1858 L=500e-9 W=3e-6
m2 net19 bl 0 0 N258 L=500e-9 W=3e-6
.ends SAVM258

.subckt SAVM259 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1859 L=500e-9 W=3e-6
m2 net19 bl 0 0 N259 L=500e-9 W=3e-6
.ends SAVM259

.subckt SAVM260 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1860 L=500e-9 W=3e-6
m2 net19 bl 0 0 N260 L=500e-9 W=3e-6
.ends SAVM260

.subckt SAVM261 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1861 L=500e-9 W=3e-6
m2 net19 bl 0 0 N261 L=500e-9 W=3e-6
.ends SAVM261

.subckt SAVM262 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1862 L=500e-9 W=3e-6
m2 net19 bl 0 0 N262 L=500e-9 W=3e-6
.ends SAVM262

.subckt SAVM263 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1863 L=500e-9 W=3e-6
m2 net19 bl 0 0 N263 L=500e-9 W=3e-6
.ends SAVM263

.subckt SAVM264 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1864 L=500e-9 W=3e-6
m2 net19 bl 0 0 N264 L=500e-9 W=3e-6
.ends SAVM264

.subckt SAVM265 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1865 L=500e-9 W=3e-6
m2 net19 bl 0 0 N265 L=500e-9 W=3e-6
.ends SAVM265

.subckt SAVM266 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1866 L=500e-9 W=3e-6
m2 net19 bl 0 0 N266 L=500e-9 W=3e-6
.ends SAVM266

.subckt SAVM267 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1867 L=500e-9 W=3e-6
m2 net19 bl 0 0 N267 L=500e-9 W=3e-6
.ends SAVM267

.subckt SAVM268 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1868 L=500e-9 W=3e-6
m2 net19 bl 0 0 N268 L=500e-9 W=3e-6
.ends SAVM268

.subckt SAVM269 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1869 L=500e-9 W=3e-6
m2 net19 bl 0 0 N269 L=500e-9 W=3e-6
.ends SAVM269

.subckt SAVM270 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1870 L=500e-9 W=3e-6
m2 net19 bl 0 0 N270 L=500e-9 W=3e-6
.ends SAVM270

.subckt SAVM271 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1871 L=500e-9 W=3e-6
m2 net19 bl 0 0 N271 L=500e-9 W=3e-6
.ends SAVM271

.subckt SAVM272 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1872 L=500e-9 W=3e-6
m2 net19 bl 0 0 N272 L=500e-9 W=3e-6
.ends SAVM272

.subckt SAVM273 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1873 L=500e-9 W=3e-6
m2 net19 bl 0 0 N273 L=500e-9 W=3e-6
.ends SAVM273

.subckt SAVM274 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1874 L=500e-9 W=3e-6
m2 net19 bl 0 0 N274 L=500e-9 W=3e-6
.ends SAVM274

.subckt SAVM275 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1875 L=500e-9 W=3e-6
m2 net19 bl 0 0 N275 L=500e-9 W=3e-6
.ends SAVM275

.subckt SAVM276 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1876 L=500e-9 W=3e-6
m2 net19 bl 0 0 N276 L=500e-9 W=3e-6
.ends SAVM276

.subckt SAVM277 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1877 L=500e-9 W=3e-6
m2 net19 bl 0 0 N277 L=500e-9 W=3e-6
.ends SAVM277

.subckt SAVM278 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1878 L=500e-9 W=3e-6
m2 net19 bl 0 0 N278 L=500e-9 W=3e-6
.ends SAVM278

.subckt SAVM279 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1879 L=500e-9 W=3e-6
m2 net19 bl 0 0 N279 L=500e-9 W=3e-6
.ends SAVM279

.subckt SAVM280 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1880 L=500e-9 W=3e-6
m2 net19 bl 0 0 N280 L=500e-9 W=3e-6
.ends SAVM280

.subckt SAVM281 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1881 L=500e-9 W=3e-6
m2 net19 bl 0 0 N281 L=500e-9 W=3e-6
.ends SAVM281

.subckt SAVM282 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1882 L=500e-9 W=3e-6
m2 net19 bl 0 0 N282 L=500e-9 W=3e-6
.ends SAVM282

.subckt SAVM283 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1883 L=500e-9 W=3e-6
m2 net19 bl 0 0 N283 L=500e-9 W=3e-6
.ends SAVM283

.subckt SAVM284 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1884 L=500e-9 W=3e-6
m2 net19 bl 0 0 N284 L=500e-9 W=3e-6
.ends SAVM284

.subckt SAVM285 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1885 L=500e-9 W=3e-6
m2 net19 bl 0 0 N285 L=500e-9 W=3e-6
.ends SAVM285

.subckt SAVM286 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1886 L=500e-9 W=3e-6
m2 net19 bl 0 0 N286 L=500e-9 W=3e-6
.ends SAVM286

.subckt SAVM287 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1887 L=500e-9 W=3e-6
m2 net19 bl 0 0 N287 L=500e-9 W=3e-6
.ends SAVM287

.subckt SAVM288 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1888 L=500e-9 W=3e-6
m2 net19 bl 0 0 N288 L=500e-9 W=3e-6
.ends SAVM288

.subckt SAVM289 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1889 L=500e-9 W=3e-6
m2 net19 bl 0 0 N289 L=500e-9 W=3e-6
.ends SAVM289

.subckt SAVM290 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1890 L=500e-9 W=3e-6
m2 net19 bl 0 0 N290 L=500e-9 W=3e-6
.ends SAVM290

.subckt SAVM291 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1891 L=500e-9 W=3e-6
m2 net19 bl 0 0 N291 L=500e-9 W=3e-6
.ends SAVM291

.subckt SAVM292 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1892 L=500e-9 W=3e-6
m2 net19 bl 0 0 N292 L=500e-9 W=3e-6
.ends SAVM292

.subckt SAVM293 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1893 L=500e-9 W=3e-6
m2 net19 bl 0 0 N293 L=500e-9 W=3e-6
.ends SAVM293

.subckt SAVM294 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1894 L=500e-9 W=3e-6
m2 net19 bl 0 0 N294 L=500e-9 W=3e-6
.ends SAVM294

.subckt SAVM295 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1895 L=500e-9 W=3e-6
m2 net19 bl 0 0 N295 L=500e-9 W=3e-6
.ends SAVM295

.subckt SAVM296 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1896 L=500e-9 W=3e-6
m2 net19 bl 0 0 N296 L=500e-9 W=3e-6
.ends SAVM296

.subckt SAVM297 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1897 L=500e-9 W=3e-6
m2 net19 bl 0 0 N297 L=500e-9 W=3e-6
.ends SAVM297

.subckt SAVM298 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1898 L=500e-9 W=3e-6
m2 net19 bl 0 0 N298 L=500e-9 W=3e-6
.ends SAVM298

.subckt SAVM299 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1899 L=500e-9 W=3e-6
m2 net19 bl 0 0 N299 L=500e-9 W=3e-6
.ends SAVM299

.subckt SAVM300 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1900 L=500e-9 W=3e-6
m2 net19 bl 0 0 N300 L=500e-9 W=3e-6
.ends SAVM300

.subckt SAVM301 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1901 L=500e-9 W=3e-6
m2 net19 bl 0 0 N301 L=500e-9 W=3e-6
.ends SAVM301

.subckt SAVM302 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1902 L=500e-9 W=3e-6
m2 net19 bl 0 0 N302 L=500e-9 W=3e-6
.ends SAVM302

.subckt SAVM303 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1903 L=500e-9 W=3e-6
m2 net19 bl 0 0 N303 L=500e-9 W=3e-6
.ends SAVM303

.subckt SAVM304 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1904 L=500e-9 W=3e-6
m2 net19 bl 0 0 N304 L=500e-9 W=3e-6
.ends SAVM304

.subckt SAVM305 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1905 L=500e-9 W=3e-6
m2 net19 bl 0 0 N305 L=500e-9 W=3e-6
.ends SAVM305

.subckt SAVM306 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1906 L=500e-9 W=3e-6
m2 net19 bl 0 0 N306 L=500e-9 W=3e-6
.ends SAVM306

.subckt SAVM307 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1907 L=500e-9 W=3e-6
m2 net19 bl 0 0 N307 L=500e-9 W=3e-6
.ends SAVM307

.subckt SAVM308 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1908 L=500e-9 W=3e-6
m2 net19 bl 0 0 N308 L=500e-9 W=3e-6
.ends SAVM308

.subckt SAVM309 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1909 L=500e-9 W=3e-6
m2 net19 bl 0 0 N309 L=500e-9 W=3e-6
.ends SAVM309

.subckt SAVM310 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1910 L=500e-9 W=3e-6
m2 net19 bl 0 0 N310 L=500e-9 W=3e-6
.ends SAVM310

.subckt SAVM311 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1911 L=500e-9 W=3e-6
m2 net19 bl 0 0 N311 L=500e-9 W=3e-6
.ends SAVM311

.subckt SAVM312 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1912 L=500e-9 W=3e-6
m2 net19 bl 0 0 N312 L=500e-9 W=3e-6
.ends SAVM312

.subckt SAVM313 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1913 L=500e-9 W=3e-6
m2 net19 bl 0 0 N313 L=500e-9 W=3e-6
.ends SAVM313

.subckt SAVM314 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1914 L=500e-9 W=3e-6
m2 net19 bl 0 0 N314 L=500e-9 W=3e-6
.ends SAVM314

.subckt SAVM315 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1915 L=500e-9 W=3e-6
m2 net19 bl 0 0 N315 L=500e-9 W=3e-6
.ends SAVM315

.subckt SAVM316 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1916 L=500e-9 W=3e-6
m2 net19 bl 0 0 N316 L=500e-9 W=3e-6
.ends SAVM316

.subckt SAVM317 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1917 L=500e-9 W=3e-6
m2 net19 bl 0 0 N317 L=500e-9 W=3e-6
.ends SAVM317

.subckt SAVM318 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1918 L=500e-9 W=3e-6
m2 net19 bl 0 0 N318 L=500e-9 W=3e-6
.ends SAVM318

.subckt SAVM319 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1919 L=500e-9 W=3e-6
m2 net19 bl 0 0 N319 L=500e-9 W=3e-6
.ends SAVM319

.subckt SAVM320 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1920 L=500e-9 W=3e-6
m2 net19 bl 0 0 N320 L=500e-9 W=3e-6
.ends SAVM320

.subckt SAVM321 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1921 L=500e-9 W=3e-6
m2 net19 bl 0 0 N321 L=500e-9 W=3e-6
.ends SAVM321

.subckt SAVM322 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1922 L=500e-9 W=3e-6
m2 net19 bl 0 0 N322 L=500e-9 W=3e-6
.ends SAVM322

.subckt SAVM323 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1923 L=500e-9 W=3e-6
m2 net19 bl 0 0 N323 L=500e-9 W=3e-6
.ends SAVM323

.subckt SAVM324 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1924 L=500e-9 W=3e-6
m2 net19 bl 0 0 N324 L=500e-9 W=3e-6
.ends SAVM324

.subckt SAVM325 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1925 L=500e-9 W=3e-6
m2 net19 bl 0 0 N325 L=500e-9 W=3e-6
.ends SAVM325

.subckt SAVM326 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1926 L=500e-9 W=3e-6
m2 net19 bl 0 0 N326 L=500e-9 W=3e-6
.ends SAVM326

.subckt SAVM327 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1927 L=500e-9 W=3e-6
m2 net19 bl 0 0 N327 L=500e-9 W=3e-6
.ends SAVM327

.subckt SAVM328 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1928 L=500e-9 W=3e-6
m2 net19 bl 0 0 N328 L=500e-9 W=3e-6
.ends SAVM328

.subckt SAVM329 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1929 L=500e-9 W=3e-6
m2 net19 bl 0 0 N329 L=500e-9 W=3e-6
.ends SAVM329

.subckt SAVM330 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1930 L=500e-9 W=3e-6
m2 net19 bl 0 0 N330 L=500e-9 W=3e-6
.ends SAVM330

.subckt SAVM331 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1931 L=500e-9 W=3e-6
m2 net19 bl 0 0 N331 L=500e-9 W=3e-6
.ends SAVM331

.subckt SAVM332 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1932 L=500e-9 W=3e-6
m2 net19 bl 0 0 N332 L=500e-9 W=3e-6
.ends SAVM332

.subckt SAVM333 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1933 L=500e-9 W=3e-6
m2 net19 bl 0 0 N333 L=500e-9 W=3e-6
.ends SAVM333

.subckt SAVM334 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1934 L=500e-9 W=3e-6
m2 net19 bl 0 0 N334 L=500e-9 W=3e-6
.ends SAVM334

.subckt SAVM335 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1935 L=500e-9 W=3e-6
m2 net19 bl 0 0 N335 L=500e-9 W=3e-6
.ends SAVM335

.subckt SAVM336 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1936 L=500e-9 W=3e-6
m2 net19 bl 0 0 N336 L=500e-9 W=3e-6
.ends SAVM336

.subckt SAVM337 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1937 L=500e-9 W=3e-6
m2 net19 bl 0 0 N337 L=500e-9 W=3e-6
.ends SAVM337

.subckt SAVM338 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1938 L=500e-9 W=3e-6
m2 net19 bl 0 0 N338 L=500e-9 W=3e-6
.ends SAVM338

.subckt SAVM339 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1939 L=500e-9 W=3e-6
m2 net19 bl 0 0 N339 L=500e-9 W=3e-6
.ends SAVM339

.subckt SAVM340 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1940 L=500e-9 W=3e-6
m2 net19 bl 0 0 N340 L=500e-9 W=3e-6
.ends SAVM340

.subckt SAVM341 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1941 L=500e-9 W=3e-6
m2 net19 bl 0 0 N341 L=500e-9 W=3e-6
.ends SAVM341

.subckt SAVM342 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1942 L=500e-9 W=3e-6
m2 net19 bl 0 0 N342 L=500e-9 W=3e-6
.ends SAVM342

.subckt SAVM343 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1943 L=500e-9 W=3e-6
m2 net19 bl 0 0 N343 L=500e-9 W=3e-6
.ends SAVM343

.subckt SAVM344 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1944 L=500e-9 W=3e-6
m2 net19 bl 0 0 N344 L=500e-9 W=3e-6
.ends SAVM344

.subckt SAVM345 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1945 L=500e-9 W=3e-6
m2 net19 bl 0 0 N345 L=500e-9 W=3e-6
.ends SAVM345

.subckt SAVM346 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1946 L=500e-9 W=3e-6
m2 net19 bl 0 0 N346 L=500e-9 W=3e-6
.ends SAVM346

.subckt SAVM347 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1947 L=500e-9 W=3e-6
m2 net19 bl 0 0 N347 L=500e-9 W=3e-6
.ends SAVM347

.subckt SAVM348 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1948 L=500e-9 W=3e-6
m2 net19 bl 0 0 N348 L=500e-9 W=3e-6
.ends SAVM348

.subckt SAVM349 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1949 L=500e-9 W=3e-6
m2 net19 bl 0 0 N349 L=500e-9 W=3e-6
.ends SAVM349

.subckt SAVM350 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1950 L=500e-9 W=3e-6
m2 net19 bl 0 0 N350 L=500e-9 W=3e-6
.ends SAVM350

.subckt SAVM351 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1951 L=500e-9 W=3e-6
m2 net19 bl 0 0 N351 L=500e-9 W=3e-6
.ends SAVM351

.subckt SAVM352 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1952 L=500e-9 W=3e-6
m2 net19 bl 0 0 N352 L=500e-9 W=3e-6
.ends SAVM352

.subckt SAVM353 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1953 L=500e-9 W=3e-6
m2 net19 bl 0 0 N353 L=500e-9 W=3e-6
.ends SAVM353

.subckt SAVM354 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1954 L=500e-9 W=3e-6
m2 net19 bl 0 0 N354 L=500e-9 W=3e-6
.ends SAVM354

.subckt SAVM355 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1955 L=500e-9 W=3e-6
m2 net19 bl 0 0 N355 L=500e-9 W=3e-6
.ends SAVM355

.subckt SAVM356 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1956 L=500e-9 W=3e-6
m2 net19 bl 0 0 N356 L=500e-9 W=3e-6
.ends SAVM356

.subckt SAVM357 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1957 L=500e-9 W=3e-6
m2 net19 bl 0 0 N357 L=500e-9 W=3e-6
.ends SAVM357

.subckt SAVM358 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1958 L=500e-9 W=3e-6
m2 net19 bl 0 0 N358 L=500e-9 W=3e-6
.ends SAVM358

.subckt SAVM359 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1959 L=500e-9 W=3e-6
m2 net19 bl 0 0 N359 L=500e-9 W=3e-6
.ends SAVM359

.subckt SAVM360 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1960 L=500e-9 W=3e-6
m2 net19 bl 0 0 N360 L=500e-9 W=3e-6
.ends SAVM360

.subckt SAVM361 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1961 L=500e-9 W=3e-6
m2 net19 bl 0 0 N361 L=500e-9 W=3e-6
.ends SAVM361

.subckt SAVM362 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1962 L=500e-9 W=3e-6
m2 net19 bl 0 0 N362 L=500e-9 W=3e-6
.ends SAVM362

.subckt SAVM363 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1963 L=500e-9 W=3e-6
m2 net19 bl 0 0 N363 L=500e-9 W=3e-6
.ends SAVM363

.subckt SAVM364 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1964 L=500e-9 W=3e-6
m2 net19 bl 0 0 N364 L=500e-9 W=3e-6
.ends SAVM364

.subckt SAVM365 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1965 L=500e-9 W=3e-6
m2 net19 bl 0 0 N365 L=500e-9 W=3e-6
.ends SAVM365

.subckt SAVM366 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1966 L=500e-9 W=3e-6
m2 net19 bl 0 0 N366 L=500e-9 W=3e-6
.ends SAVM366

.subckt SAVM367 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1967 L=500e-9 W=3e-6
m2 net19 bl 0 0 N367 L=500e-9 W=3e-6
.ends SAVM367

.subckt SAVM368 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1968 L=500e-9 W=3e-6
m2 net19 bl 0 0 N368 L=500e-9 W=3e-6
.ends SAVM368

.subckt SAVM369 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1969 L=500e-9 W=3e-6
m2 net19 bl 0 0 N369 L=500e-9 W=3e-6
.ends SAVM369

.subckt SAVM370 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1970 L=500e-9 W=3e-6
m2 net19 bl 0 0 N370 L=500e-9 W=3e-6
.ends SAVM370

.subckt SAVM371 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1971 L=500e-9 W=3e-6
m2 net19 bl 0 0 N371 L=500e-9 W=3e-6
.ends SAVM371

.subckt SAVM372 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1972 L=500e-9 W=3e-6
m2 net19 bl 0 0 N372 L=500e-9 W=3e-6
.ends SAVM372

.subckt SAVM373 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1973 L=500e-9 W=3e-6
m2 net19 bl 0 0 N373 L=500e-9 W=3e-6
.ends SAVM373

.subckt SAVM374 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1974 L=500e-9 W=3e-6
m2 net19 bl 0 0 N374 L=500e-9 W=3e-6
.ends SAVM374

.subckt SAVM375 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1975 L=500e-9 W=3e-6
m2 net19 bl 0 0 N375 L=500e-9 W=3e-6
.ends SAVM375

.subckt SAVM376 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1976 L=500e-9 W=3e-6
m2 net19 bl 0 0 N376 L=500e-9 W=3e-6
.ends SAVM376

.subckt SAVM377 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1977 L=500e-9 W=3e-6
m2 net19 bl 0 0 N377 L=500e-9 W=3e-6
.ends SAVM377

.subckt SAVM378 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1978 L=500e-9 W=3e-6
m2 net19 bl 0 0 N378 L=500e-9 W=3e-6
.ends SAVM378

.subckt SAVM379 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1979 L=500e-9 W=3e-6
m2 net19 bl 0 0 N379 L=500e-9 W=3e-6
.ends SAVM379

.subckt SAVM380 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1980 L=500e-9 W=3e-6
m2 net19 bl 0 0 N380 L=500e-9 W=3e-6
.ends SAVM380

.subckt SAVM381 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1981 L=500e-9 W=3e-6
m2 net19 bl 0 0 N381 L=500e-9 W=3e-6
.ends SAVM381

.subckt SAVM382 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1982 L=500e-9 W=3e-6
m2 net19 bl 0 0 N382 L=500e-9 W=3e-6
.ends SAVM382

.subckt SAVM383 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1983 L=500e-9 W=3e-6
m2 net19 bl 0 0 N383 L=500e-9 W=3e-6
.ends SAVM383

.subckt SAVM384 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1984 L=500e-9 W=3e-6
m2 net19 bl 0 0 N384 L=500e-9 W=3e-6
.ends SAVM384

.subckt SAVM385 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1985 L=500e-9 W=3e-6
m2 net19 bl 0 0 N385 L=500e-9 W=3e-6
.ends SAVM385

.subckt SAVM386 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1986 L=500e-9 W=3e-6
m2 net19 bl 0 0 N386 L=500e-9 W=3e-6
.ends SAVM386

.subckt SAVM387 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1987 L=500e-9 W=3e-6
m2 net19 bl 0 0 N387 L=500e-9 W=3e-6
.ends SAVM387

.subckt SAVM388 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1988 L=500e-9 W=3e-6
m2 net19 bl 0 0 N388 L=500e-9 W=3e-6
.ends SAVM388

.subckt SAVM389 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1989 L=500e-9 W=3e-6
m2 net19 bl 0 0 N389 L=500e-9 W=3e-6
.ends SAVM389

.subckt SAVM390 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1990 L=500e-9 W=3e-6
m2 net19 bl 0 0 N390 L=500e-9 W=3e-6
.ends SAVM390

.subckt SAVM391 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1991 L=500e-9 W=3e-6
m2 net19 bl 0 0 N391 L=500e-9 W=3e-6
.ends SAVM391

.subckt SAVM392 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1992 L=500e-9 W=3e-6
m2 net19 bl 0 0 N392 L=500e-9 W=3e-6
.ends SAVM392

.subckt SAVM393 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1993 L=500e-9 W=3e-6
m2 net19 bl 0 0 N393 L=500e-9 W=3e-6
.ends SAVM393

.subckt SAVM394 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1994 L=500e-9 W=3e-6
m2 net19 bl 0 0 N394 L=500e-9 W=3e-6
.ends SAVM394

.subckt SAVM395 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1995 L=500e-9 W=3e-6
m2 net19 bl 0 0 N395 L=500e-9 W=3e-6
.ends SAVM395

.subckt SAVM396 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1996 L=500e-9 W=3e-6
m2 net19 bl 0 0 N396 L=500e-9 W=3e-6
.ends SAVM396

.subckt SAVM397 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1997 L=500e-9 W=3e-6
m2 net19 bl 0 0 N397 L=500e-9 W=3e-6
.ends SAVM397

.subckt SAVM398 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1998 L=500e-9 W=3e-6
m2 net19 bl 0 0 N398 L=500e-9 W=3e-6
.ends SAVM398

.subckt SAVM399 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N1999 L=500e-9 W=3e-6
m2 net19 bl 0 0 N399 L=500e-9 W=3e-6
.ends SAVM399

.subckt SAVM400 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2000 L=500e-9 W=3e-6
m2 net19 bl 0 0 N400 L=500e-9 W=3e-6
.ends SAVM400

.subckt SAVM401 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2001 L=500e-9 W=3e-6
m2 net19 bl 0 0 N401 L=500e-9 W=3e-6
.ends SAVM401

.subckt SAVM402 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2002 L=500e-9 W=3e-6
m2 net19 bl 0 0 N402 L=500e-9 W=3e-6
.ends SAVM402

.subckt SAVM403 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2003 L=500e-9 W=3e-6
m2 net19 bl 0 0 N403 L=500e-9 W=3e-6
.ends SAVM403

.subckt SAVM404 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2004 L=500e-9 W=3e-6
m2 net19 bl 0 0 N404 L=500e-9 W=3e-6
.ends SAVM404

.subckt SAVM405 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2005 L=500e-9 W=3e-6
m2 net19 bl 0 0 N405 L=500e-9 W=3e-6
.ends SAVM405

.subckt SAVM406 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2006 L=500e-9 W=3e-6
m2 net19 bl 0 0 N406 L=500e-9 W=3e-6
.ends SAVM406

.subckt SAVM407 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2007 L=500e-9 W=3e-6
m2 net19 bl 0 0 N407 L=500e-9 W=3e-6
.ends SAVM407

.subckt SAVM408 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2008 L=500e-9 W=3e-6
m2 net19 bl 0 0 N408 L=500e-9 W=3e-6
.ends SAVM408

.subckt SAVM409 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2009 L=500e-9 W=3e-6
m2 net19 bl 0 0 N409 L=500e-9 W=3e-6
.ends SAVM409

.subckt SAVM410 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2010 L=500e-9 W=3e-6
m2 net19 bl 0 0 N410 L=500e-9 W=3e-6
.ends SAVM410

.subckt SAVM411 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2011 L=500e-9 W=3e-6
m2 net19 bl 0 0 N411 L=500e-9 W=3e-6
.ends SAVM411

.subckt SAVM412 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2012 L=500e-9 W=3e-6
m2 net19 bl 0 0 N412 L=500e-9 W=3e-6
.ends SAVM412

.subckt SAVM413 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2013 L=500e-9 W=3e-6
m2 net19 bl 0 0 N413 L=500e-9 W=3e-6
.ends SAVM413

.subckt SAVM414 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2014 L=500e-9 W=3e-6
m2 net19 bl 0 0 N414 L=500e-9 W=3e-6
.ends SAVM414

.subckt SAVM415 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2015 L=500e-9 W=3e-6
m2 net19 bl 0 0 N415 L=500e-9 W=3e-6
.ends SAVM415

.subckt SAVM416 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2016 L=500e-9 W=3e-6
m2 net19 bl 0 0 N416 L=500e-9 W=3e-6
.ends SAVM416

.subckt SAVM417 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2017 L=500e-9 W=3e-6
m2 net19 bl 0 0 N417 L=500e-9 W=3e-6
.ends SAVM417

.subckt SAVM418 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2018 L=500e-9 W=3e-6
m2 net19 bl 0 0 N418 L=500e-9 W=3e-6
.ends SAVM418

.subckt SAVM419 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2019 L=500e-9 W=3e-6
m2 net19 bl 0 0 N419 L=500e-9 W=3e-6
.ends SAVM419

.subckt SAVM420 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2020 L=500e-9 W=3e-6
m2 net19 bl 0 0 N420 L=500e-9 W=3e-6
.ends SAVM420

.subckt SAVM421 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2021 L=500e-9 W=3e-6
m2 net19 bl 0 0 N421 L=500e-9 W=3e-6
.ends SAVM421

.subckt SAVM422 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2022 L=500e-9 W=3e-6
m2 net19 bl 0 0 N422 L=500e-9 W=3e-6
.ends SAVM422

.subckt SAVM423 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2023 L=500e-9 W=3e-6
m2 net19 bl 0 0 N423 L=500e-9 W=3e-6
.ends SAVM423

.subckt SAVM424 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2024 L=500e-9 W=3e-6
m2 net19 bl 0 0 N424 L=500e-9 W=3e-6
.ends SAVM424

.subckt SAVM425 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2025 L=500e-9 W=3e-6
m2 net19 bl 0 0 N425 L=500e-9 W=3e-6
.ends SAVM425

.subckt SAVM426 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2026 L=500e-9 W=3e-6
m2 net19 bl 0 0 N426 L=500e-9 W=3e-6
.ends SAVM426

.subckt SAVM427 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2027 L=500e-9 W=3e-6
m2 net19 bl 0 0 N427 L=500e-9 W=3e-6
.ends SAVM427

.subckt SAVM428 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2028 L=500e-9 W=3e-6
m2 net19 bl 0 0 N428 L=500e-9 W=3e-6
.ends SAVM428

.subckt SAVM429 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2029 L=500e-9 W=3e-6
m2 net19 bl 0 0 N429 L=500e-9 W=3e-6
.ends SAVM429

.subckt SAVM430 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2030 L=500e-9 W=3e-6
m2 net19 bl 0 0 N430 L=500e-9 W=3e-6
.ends SAVM430

.subckt SAVM431 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2031 L=500e-9 W=3e-6
m2 net19 bl 0 0 N431 L=500e-9 W=3e-6
.ends SAVM431

.subckt SAVM432 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2032 L=500e-9 W=3e-6
m2 net19 bl 0 0 N432 L=500e-9 W=3e-6
.ends SAVM432

.subckt SAVM433 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2033 L=500e-9 W=3e-6
m2 net19 bl 0 0 N433 L=500e-9 W=3e-6
.ends SAVM433

.subckt SAVM434 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2034 L=500e-9 W=3e-6
m2 net19 bl 0 0 N434 L=500e-9 W=3e-6
.ends SAVM434

.subckt SAVM435 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2035 L=500e-9 W=3e-6
m2 net19 bl 0 0 N435 L=500e-9 W=3e-6
.ends SAVM435

.subckt SAVM436 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2036 L=500e-9 W=3e-6
m2 net19 bl 0 0 N436 L=500e-9 W=3e-6
.ends SAVM436

.subckt SAVM437 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2037 L=500e-9 W=3e-6
m2 net19 bl 0 0 N437 L=500e-9 W=3e-6
.ends SAVM437

.subckt SAVM438 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2038 L=500e-9 W=3e-6
m2 net19 bl 0 0 N438 L=500e-9 W=3e-6
.ends SAVM438

.subckt SAVM439 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2039 L=500e-9 W=3e-6
m2 net19 bl 0 0 N439 L=500e-9 W=3e-6
.ends SAVM439

.subckt SAVM440 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2040 L=500e-9 W=3e-6
m2 net19 bl 0 0 N440 L=500e-9 W=3e-6
.ends SAVM440

.subckt SAVM441 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2041 L=500e-9 W=3e-6
m2 net19 bl 0 0 N441 L=500e-9 W=3e-6
.ends SAVM441

.subckt SAVM442 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2042 L=500e-9 W=3e-6
m2 net19 bl 0 0 N442 L=500e-9 W=3e-6
.ends SAVM442

.subckt SAVM443 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2043 L=500e-9 W=3e-6
m2 net19 bl 0 0 N443 L=500e-9 W=3e-6
.ends SAVM443

.subckt SAVM444 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2044 L=500e-9 W=3e-6
m2 net19 bl 0 0 N444 L=500e-9 W=3e-6
.ends SAVM444

.subckt SAVM445 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2045 L=500e-9 W=3e-6
m2 net19 bl 0 0 N445 L=500e-9 W=3e-6
.ends SAVM445

.subckt SAVM446 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2046 L=500e-9 W=3e-6
m2 net19 bl 0 0 N446 L=500e-9 W=3e-6
.ends SAVM446

.subckt SAVM447 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2047 L=500e-9 W=3e-6
m2 net19 bl 0 0 N447 L=500e-9 W=3e-6
.ends SAVM447

.subckt SAVM448 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2048 L=500e-9 W=3e-6
m2 net19 bl 0 0 N448 L=500e-9 W=3e-6
.ends SAVM448

.subckt SAVM449 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2049 L=500e-9 W=3e-6
m2 net19 bl 0 0 N449 L=500e-9 W=3e-6
.ends SAVM449

.subckt SAVM450 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2050 L=500e-9 W=3e-6
m2 net19 bl 0 0 N450 L=500e-9 W=3e-6
.ends SAVM450

.subckt SAVM451 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2051 L=500e-9 W=3e-6
m2 net19 bl 0 0 N451 L=500e-9 W=3e-6
.ends SAVM451

.subckt SAVM452 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2052 L=500e-9 W=3e-6
m2 net19 bl 0 0 N452 L=500e-9 W=3e-6
.ends SAVM452

.subckt SAVM453 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2053 L=500e-9 W=3e-6
m2 net19 bl 0 0 N453 L=500e-9 W=3e-6
.ends SAVM453

.subckt SAVM454 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2054 L=500e-9 W=3e-6
m2 net19 bl 0 0 N454 L=500e-9 W=3e-6
.ends SAVM454

.subckt SAVM455 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2055 L=500e-9 W=3e-6
m2 net19 bl 0 0 N455 L=500e-9 W=3e-6
.ends SAVM455

.subckt SAVM456 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2056 L=500e-9 W=3e-6
m2 net19 bl 0 0 N456 L=500e-9 W=3e-6
.ends SAVM456

.subckt SAVM457 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2057 L=500e-9 W=3e-6
m2 net19 bl 0 0 N457 L=500e-9 W=3e-6
.ends SAVM457

.subckt SAVM458 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2058 L=500e-9 W=3e-6
m2 net19 bl 0 0 N458 L=500e-9 W=3e-6
.ends SAVM458

.subckt SAVM459 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2059 L=500e-9 W=3e-6
m2 net19 bl 0 0 N459 L=500e-9 W=3e-6
.ends SAVM459

.subckt SAVM460 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2060 L=500e-9 W=3e-6
m2 net19 bl 0 0 N460 L=500e-9 W=3e-6
.ends SAVM460

.subckt SAVM461 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2061 L=500e-9 W=3e-6
m2 net19 bl 0 0 N461 L=500e-9 W=3e-6
.ends SAVM461

.subckt SAVM462 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2062 L=500e-9 W=3e-6
m2 net19 bl 0 0 N462 L=500e-9 W=3e-6
.ends SAVM462

.subckt SAVM463 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2063 L=500e-9 W=3e-6
m2 net19 bl 0 0 N463 L=500e-9 W=3e-6
.ends SAVM463

.subckt SAVM464 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2064 L=500e-9 W=3e-6
m2 net19 bl 0 0 N464 L=500e-9 W=3e-6
.ends SAVM464

.subckt SAVM465 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2065 L=500e-9 W=3e-6
m2 net19 bl 0 0 N465 L=500e-9 W=3e-6
.ends SAVM465

.subckt SAVM466 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2066 L=500e-9 W=3e-6
m2 net19 bl 0 0 N466 L=500e-9 W=3e-6
.ends SAVM466

.subckt SAVM467 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2067 L=500e-9 W=3e-6
m2 net19 bl 0 0 N467 L=500e-9 W=3e-6
.ends SAVM467

.subckt SAVM468 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2068 L=500e-9 W=3e-6
m2 net19 bl 0 0 N468 L=500e-9 W=3e-6
.ends SAVM468

.subckt SAVM469 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2069 L=500e-9 W=3e-6
m2 net19 bl 0 0 N469 L=500e-9 W=3e-6
.ends SAVM469

.subckt SAVM470 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2070 L=500e-9 W=3e-6
m2 net19 bl 0 0 N470 L=500e-9 W=3e-6
.ends SAVM470

.subckt SAVM471 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2071 L=500e-9 W=3e-6
m2 net19 bl 0 0 N471 L=500e-9 W=3e-6
.ends SAVM471

.subckt SAVM472 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2072 L=500e-9 W=3e-6
m2 net19 bl 0 0 N472 L=500e-9 W=3e-6
.ends SAVM472

.subckt SAVM473 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2073 L=500e-9 W=3e-6
m2 net19 bl 0 0 N473 L=500e-9 W=3e-6
.ends SAVM473

.subckt SAVM474 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2074 L=500e-9 W=3e-6
m2 net19 bl 0 0 N474 L=500e-9 W=3e-6
.ends SAVM474

.subckt SAVM475 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2075 L=500e-9 W=3e-6
m2 net19 bl 0 0 N475 L=500e-9 W=3e-6
.ends SAVM475

.subckt SAVM476 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2076 L=500e-9 W=3e-6
m2 net19 bl 0 0 N476 L=500e-9 W=3e-6
.ends SAVM476

.subckt SAVM477 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2077 L=500e-9 W=3e-6
m2 net19 bl 0 0 N477 L=500e-9 W=3e-6
.ends SAVM477

.subckt SAVM478 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2078 L=500e-9 W=3e-6
m2 net19 bl 0 0 N478 L=500e-9 W=3e-6
.ends SAVM478

.subckt SAVM479 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2079 L=500e-9 W=3e-6
m2 net19 bl 0 0 N479 L=500e-9 W=3e-6
.ends SAVM479

.subckt SAVM480 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2080 L=500e-9 W=3e-6
m2 net19 bl 0 0 N480 L=500e-9 W=3e-6
.ends SAVM480

.subckt SAVM481 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2081 L=500e-9 W=3e-6
m2 net19 bl 0 0 N481 L=500e-9 W=3e-6
.ends SAVM481

.subckt SAVM482 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2082 L=500e-9 W=3e-6
m2 net19 bl 0 0 N482 L=500e-9 W=3e-6
.ends SAVM482

.subckt SAVM483 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2083 L=500e-9 W=3e-6
m2 net19 bl 0 0 N483 L=500e-9 W=3e-6
.ends SAVM483

.subckt SAVM484 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2084 L=500e-9 W=3e-6
m2 net19 bl 0 0 N484 L=500e-9 W=3e-6
.ends SAVM484

.subckt SAVM485 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2085 L=500e-9 W=3e-6
m2 net19 bl 0 0 N485 L=500e-9 W=3e-6
.ends SAVM485

.subckt SAVM486 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2086 L=500e-9 W=3e-6
m2 net19 bl 0 0 N486 L=500e-9 W=3e-6
.ends SAVM486

.subckt SAVM487 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2087 L=500e-9 W=3e-6
m2 net19 bl 0 0 N487 L=500e-9 W=3e-6
.ends SAVM487

.subckt SAVM488 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2088 L=500e-9 W=3e-6
m2 net19 bl 0 0 N488 L=500e-9 W=3e-6
.ends SAVM488

.subckt SAVM489 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2089 L=500e-9 W=3e-6
m2 net19 bl 0 0 N489 L=500e-9 W=3e-6
.ends SAVM489

.subckt SAVM490 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2090 L=500e-9 W=3e-6
m2 net19 bl 0 0 N490 L=500e-9 W=3e-6
.ends SAVM490

.subckt SAVM491 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2091 L=500e-9 W=3e-6
m2 net19 bl 0 0 N491 L=500e-9 W=3e-6
.ends SAVM491

.subckt SAVM492 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2092 L=500e-9 W=3e-6
m2 net19 bl 0 0 N492 L=500e-9 W=3e-6
.ends SAVM492

.subckt SAVM493 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2093 L=500e-9 W=3e-6
m2 net19 bl 0 0 N493 L=500e-9 W=3e-6
.ends SAVM493

.subckt SAVM494 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2094 L=500e-9 W=3e-6
m2 net19 bl 0 0 N494 L=500e-9 W=3e-6
.ends SAVM494

.subckt SAVM495 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2095 L=500e-9 W=3e-6
m2 net19 bl 0 0 N495 L=500e-9 W=3e-6
.ends SAVM495

.subckt SAVM496 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2096 L=500e-9 W=3e-6
m2 net19 bl 0 0 N496 L=500e-9 W=3e-6
.ends SAVM496

.subckt SAVM497 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2097 L=500e-9 W=3e-6
m2 net19 bl 0 0 N497 L=500e-9 W=3e-6
.ends SAVM497

.subckt SAVM498 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2098 L=500e-9 W=3e-6
m2 net19 bl 0 0 N498 L=500e-9 W=3e-6
.ends SAVM498

.subckt SAVM499 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2099 L=500e-9 W=3e-6
m2 net19 bl 0 0 N499 L=500e-9 W=3e-6
.ends SAVM499

.subckt SAVM500 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2100 L=500e-9 W=3e-6
m2 net19 bl 0 0 N500 L=500e-9 W=3e-6
.ends SAVM500

.subckt SAVM501 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2101 L=500e-9 W=3e-6
m2 net19 bl 0 0 N501 L=500e-9 W=3e-6
.ends SAVM501

.subckt SAVM502 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2102 L=500e-9 W=3e-6
m2 net19 bl 0 0 N502 L=500e-9 W=3e-6
.ends SAVM502

.subckt SAVM503 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2103 L=500e-9 W=3e-6
m2 net19 bl 0 0 N503 L=500e-9 W=3e-6
.ends SAVM503

.subckt SAVM504 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2104 L=500e-9 W=3e-6
m2 net19 bl 0 0 N504 L=500e-9 W=3e-6
.ends SAVM504

.subckt SAVM505 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2105 L=500e-9 W=3e-6
m2 net19 bl 0 0 N505 L=500e-9 W=3e-6
.ends SAVM505

.subckt SAVM506 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2106 L=500e-9 W=3e-6
m2 net19 bl 0 0 N506 L=500e-9 W=3e-6
.ends SAVM506

.subckt SAVM507 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2107 L=500e-9 W=3e-6
m2 net19 bl 0 0 N507 L=500e-9 W=3e-6
.ends SAVM507

.subckt SAVM508 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2108 L=500e-9 W=3e-6
m2 net19 bl 0 0 N508 L=500e-9 W=3e-6
.ends SAVM508

.subckt SAVM509 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2109 L=500e-9 W=3e-6
m2 net19 bl 0 0 N509 L=500e-9 W=3e-6
.ends SAVM509

.subckt SAVM510 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2110 L=500e-9 W=3e-6
m2 net19 bl 0 0 N510 L=500e-9 W=3e-6
.ends SAVM510

.subckt SAVM511 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2111 L=500e-9 W=3e-6
m2 net19 bl 0 0 N511 L=500e-9 W=3e-6
.ends SAVM511

.subckt SAVM512 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2112 L=500e-9 W=3e-6
m2 net19 bl 0 0 N512 L=500e-9 W=3e-6
.ends SAVM512

.subckt SAVM513 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2113 L=500e-9 W=3e-6
m2 net19 bl 0 0 N513 L=500e-9 W=3e-6
.ends SAVM513

.subckt SAVM514 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2114 L=500e-9 W=3e-6
m2 net19 bl 0 0 N514 L=500e-9 W=3e-6
.ends SAVM514

.subckt SAVM515 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2115 L=500e-9 W=3e-6
m2 net19 bl 0 0 N515 L=500e-9 W=3e-6
.ends SAVM515

.subckt SAVM516 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2116 L=500e-9 W=3e-6
m2 net19 bl 0 0 N516 L=500e-9 W=3e-6
.ends SAVM516

.subckt SAVM517 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2117 L=500e-9 W=3e-6
m2 net19 bl 0 0 N517 L=500e-9 W=3e-6
.ends SAVM517

.subckt SAVM518 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2118 L=500e-9 W=3e-6
m2 net19 bl 0 0 N518 L=500e-9 W=3e-6
.ends SAVM518

.subckt SAVM519 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2119 L=500e-9 W=3e-6
m2 net19 bl 0 0 N519 L=500e-9 W=3e-6
.ends SAVM519

.subckt SAVM520 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2120 L=500e-9 W=3e-6
m2 net19 bl 0 0 N520 L=500e-9 W=3e-6
.ends SAVM520

.subckt SAVM521 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2121 L=500e-9 W=3e-6
m2 net19 bl 0 0 N521 L=500e-9 W=3e-6
.ends SAVM521

.subckt SAVM522 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2122 L=500e-9 W=3e-6
m2 net19 bl 0 0 N522 L=500e-9 W=3e-6
.ends SAVM522

.subckt SAVM523 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2123 L=500e-9 W=3e-6
m2 net19 bl 0 0 N523 L=500e-9 W=3e-6
.ends SAVM523

.subckt SAVM524 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2124 L=500e-9 W=3e-6
m2 net19 bl 0 0 N524 L=500e-9 W=3e-6
.ends SAVM524

.subckt SAVM525 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2125 L=500e-9 W=3e-6
m2 net19 bl 0 0 N525 L=500e-9 W=3e-6
.ends SAVM525

.subckt SAVM526 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2126 L=500e-9 W=3e-6
m2 net19 bl 0 0 N526 L=500e-9 W=3e-6
.ends SAVM526

.subckt SAVM527 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2127 L=500e-9 W=3e-6
m2 net19 bl 0 0 N527 L=500e-9 W=3e-6
.ends SAVM527

.subckt SAVM528 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2128 L=500e-9 W=3e-6
m2 net19 bl 0 0 N528 L=500e-9 W=3e-6
.ends SAVM528

.subckt SAVM529 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2129 L=500e-9 W=3e-6
m2 net19 bl 0 0 N529 L=500e-9 W=3e-6
.ends SAVM529

.subckt SAVM530 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2130 L=500e-9 W=3e-6
m2 net19 bl 0 0 N530 L=500e-9 W=3e-6
.ends SAVM530

.subckt SAVM531 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2131 L=500e-9 W=3e-6
m2 net19 bl 0 0 N531 L=500e-9 W=3e-6
.ends SAVM531

.subckt SAVM532 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2132 L=500e-9 W=3e-6
m2 net19 bl 0 0 N532 L=500e-9 W=3e-6
.ends SAVM532

.subckt SAVM533 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2133 L=500e-9 W=3e-6
m2 net19 bl 0 0 N533 L=500e-9 W=3e-6
.ends SAVM533

.subckt SAVM534 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2134 L=500e-9 W=3e-6
m2 net19 bl 0 0 N534 L=500e-9 W=3e-6
.ends SAVM534

.subckt SAVM535 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2135 L=500e-9 W=3e-6
m2 net19 bl 0 0 N535 L=500e-9 W=3e-6
.ends SAVM535

.subckt SAVM536 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2136 L=500e-9 W=3e-6
m2 net19 bl 0 0 N536 L=500e-9 W=3e-6
.ends SAVM536

.subckt SAVM537 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2137 L=500e-9 W=3e-6
m2 net19 bl 0 0 N537 L=500e-9 W=3e-6
.ends SAVM537

.subckt SAVM538 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2138 L=500e-9 W=3e-6
m2 net19 bl 0 0 N538 L=500e-9 W=3e-6
.ends SAVM538

.subckt SAVM539 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2139 L=500e-9 W=3e-6
m2 net19 bl 0 0 N539 L=500e-9 W=3e-6
.ends SAVM539

.subckt SAVM540 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2140 L=500e-9 W=3e-6
m2 net19 bl 0 0 N540 L=500e-9 W=3e-6
.ends SAVM540

.subckt SAVM541 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2141 L=500e-9 W=3e-6
m2 net19 bl 0 0 N541 L=500e-9 W=3e-6
.ends SAVM541

.subckt SAVM542 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2142 L=500e-9 W=3e-6
m2 net19 bl 0 0 N542 L=500e-9 W=3e-6
.ends SAVM542

.subckt SAVM543 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2143 L=500e-9 W=3e-6
m2 net19 bl 0 0 N543 L=500e-9 W=3e-6
.ends SAVM543

.subckt SAVM544 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2144 L=500e-9 W=3e-6
m2 net19 bl 0 0 N544 L=500e-9 W=3e-6
.ends SAVM544

.subckt SAVM545 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2145 L=500e-9 W=3e-6
m2 net19 bl 0 0 N545 L=500e-9 W=3e-6
.ends SAVM545

.subckt SAVM546 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2146 L=500e-9 W=3e-6
m2 net19 bl 0 0 N546 L=500e-9 W=3e-6
.ends SAVM546

.subckt SAVM547 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2147 L=500e-9 W=3e-6
m2 net19 bl 0 0 N547 L=500e-9 W=3e-6
.ends SAVM547

.subckt SAVM548 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2148 L=500e-9 W=3e-6
m2 net19 bl 0 0 N548 L=500e-9 W=3e-6
.ends SAVM548

.subckt SAVM549 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2149 L=500e-9 W=3e-6
m2 net19 bl 0 0 N549 L=500e-9 W=3e-6
.ends SAVM549

.subckt SAVM550 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2150 L=500e-9 W=3e-6
m2 net19 bl 0 0 N550 L=500e-9 W=3e-6
.ends SAVM550

.subckt SAVM551 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2151 L=500e-9 W=3e-6
m2 net19 bl 0 0 N551 L=500e-9 W=3e-6
.ends SAVM551

.subckt SAVM552 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2152 L=500e-9 W=3e-6
m2 net19 bl 0 0 N552 L=500e-9 W=3e-6
.ends SAVM552

.subckt SAVM553 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2153 L=500e-9 W=3e-6
m2 net19 bl 0 0 N553 L=500e-9 W=3e-6
.ends SAVM553

.subckt SAVM554 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2154 L=500e-9 W=3e-6
m2 net19 bl 0 0 N554 L=500e-9 W=3e-6
.ends SAVM554

.subckt SAVM555 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2155 L=500e-9 W=3e-6
m2 net19 bl 0 0 N555 L=500e-9 W=3e-6
.ends SAVM555

.subckt SAVM556 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2156 L=500e-9 W=3e-6
m2 net19 bl 0 0 N556 L=500e-9 W=3e-6
.ends SAVM556

.subckt SAVM557 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2157 L=500e-9 W=3e-6
m2 net19 bl 0 0 N557 L=500e-9 W=3e-6
.ends SAVM557

.subckt SAVM558 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2158 L=500e-9 W=3e-6
m2 net19 bl 0 0 N558 L=500e-9 W=3e-6
.ends SAVM558

.subckt SAVM559 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2159 L=500e-9 W=3e-6
m2 net19 bl 0 0 N559 L=500e-9 W=3e-6
.ends SAVM559

.subckt SAVM560 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2160 L=500e-9 W=3e-6
m2 net19 bl 0 0 N560 L=500e-9 W=3e-6
.ends SAVM560

.subckt SAVM561 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2161 L=500e-9 W=3e-6
m2 net19 bl 0 0 N561 L=500e-9 W=3e-6
.ends SAVM561

.subckt SAVM562 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2162 L=500e-9 W=3e-6
m2 net19 bl 0 0 N562 L=500e-9 W=3e-6
.ends SAVM562

.subckt SAVM563 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2163 L=500e-9 W=3e-6
m2 net19 bl 0 0 N563 L=500e-9 W=3e-6
.ends SAVM563

.subckt SAVM564 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2164 L=500e-9 W=3e-6
m2 net19 bl 0 0 N564 L=500e-9 W=3e-6
.ends SAVM564

.subckt SAVM565 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2165 L=500e-9 W=3e-6
m2 net19 bl 0 0 N565 L=500e-9 W=3e-6
.ends SAVM565

.subckt SAVM566 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2166 L=500e-9 W=3e-6
m2 net19 bl 0 0 N566 L=500e-9 W=3e-6
.ends SAVM566

.subckt SAVM567 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2167 L=500e-9 W=3e-6
m2 net19 bl 0 0 N567 L=500e-9 W=3e-6
.ends SAVM567

.subckt SAVM568 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2168 L=500e-9 W=3e-6
m2 net19 bl 0 0 N568 L=500e-9 W=3e-6
.ends SAVM568

.subckt SAVM569 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2169 L=500e-9 W=3e-6
m2 net19 bl 0 0 N569 L=500e-9 W=3e-6
.ends SAVM569

.subckt SAVM570 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2170 L=500e-9 W=3e-6
m2 net19 bl 0 0 N570 L=500e-9 W=3e-6
.ends SAVM570

.subckt SAVM571 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2171 L=500e-9 W=3e-6
m2 net19 bl 0 0 N571 L=500e-9 W=3e-6
.ends SAVM571

.subckt SAVM572 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2172 L=500e-9 W=3e-6
m2 net19 bl 0 0 N572 L=500e-9 W=3e-6
.ends SAVM572

.subckt SAVM573 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2173 L=500e-9 W=3e-6
m2 net19 bl 0 0 N573 L=500e-9 W=3e-6
.ends SAVM573

.subckt SAVM574 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2174 L=500e-9 W=3e-6
m2 net19 bl 0 0 N574 L=500e-9 W=3e-6
.ends SAVM574

.subckt SAVM575 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2175 L=500e-9 W=3e-6
m2 net19 bl 0 0 N575 L=500e-9 W=3e-6
.ends SAVM575

.subckt SAVM576 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2176 L=500e-9 W=3e-6
m2 net19 bl 0 0 N576 L=500e-9 W=3e-6
.ends SAVM576

.subckt SAVM577 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2177 L=500e-9 W=3e-6
m2 net19 bl 0 0 N577 L=500e-9 W=3e-6
.ends SAVM577

.subckt SAVM578 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2178 L=500e-9 W=3e-6
m2 net19 bl 0 0 N578 L=500e-9 W=3e-6
.ends SAVM578

.subckt SAVM579 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2179 L=500e-9 W=3e-6
m2 net19 bl 0 0 N579 L=500e-9 W=3e-6
.ends SAVM579

.subckt SAVM580 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2180 L=500e-9 W=3e-6
m2 net19 bl 0 0 N580 L=500e-9 W=3e-6
.ends SAVM580

.subckt SAVM581 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2181 L=500e-9 W=3e-6
m2 net19 bl 0 0 N581 L=500e-9 W=3e-6
.ends SAVM581

.subckt SAVM582 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2182 L=500e-9 W=3e-6
m2 net19 bl 0 0 N582 L=500e-9 W=3e-6
.ends SAVM582

.subckt SAVM583 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2183 L=500e-9 W=3e-6
m2 net19 bl 0 0 N583 L=500e-9 W=3e-6
.ends SAVM583

.subckt SAVM584 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2184 L=500e-9 W=3e-6
m2 net19 bl 0 0 N584 L=500e-9 W=3e-6
.ends SAVM584

.subckt SAVM585 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2185 L=500e-9 W=3e-6
m2 net19 bl 0 0 N585 L=500e-9 W=3e-6
.ends SAVM585

.subckt SAVM586 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2186 L=500e-9 W=3e-6
m2 net19 bl 0 0 N586 L=500e-9 W=3e-6
.ends SAVM586

.subckt SAVM587 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2187 L=500e-9 W=3e-6
m2 net19 bl 0 0 N587 L=500e-9 W=3e-6
.ends SAVM587

.subckt SAVM588 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2188 L=500e-9 W=3e-6
m2 net19 bl 0 0 N588 L=500e-9 W=3e-6
.ends SAVM588

.subckt SAVM589 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2189 L=500e-9 W=3e-6
m2 net19 bl 0 0 N589 L=500e-9 W=3e-6
.ends SAVM589

.subckt SAVM590 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2190 L=500e-9 W=3e-6
m2 net19 bl 0 0 N590 L=500e-9 W=3e-6
.ends SAVM590

.subckt SAVM591 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2191 L=500e-9 W=3e-6
m2 net19 bl 0 0 N591 L=500e-9 W=3e-6
.ends SAVM591

.subckt SAVM592 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2192 L=500e-9 W=3e-6
m2 net19 bl 0 0 N592 L=500e-9 W=3e-6
.ends SAVM592

.subckt SAVM593 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2193 L=500e-9 W=3e-6
m2 net19 bl 0 0 N593 L=500e-9 W=3e-6
.ends SAVM593

.subckt SAVM594 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2194 L=500e-9 W=3e-6
m2 net19 bl 0 0 N594 L=500e-9 W=3e-6
.ends SAVM594

.subckt SAVM595 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2195 L=500e-9 W=3e-6
m2 net19 bl 0 0 N595 L=500e-9 W=3e-6
.ends SAVM595

.subckt SAVM596 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2196 L=500e-9 W=3e-6
m2 net19 bl 0 0 N596 L=500e-9 W=3e-6
.ends SAVM596

.subckt SAVM597 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2197 L=500e-9 W=3e-6
m2 net19 bl 0 0 N597 L=500e-9 W=3e-6
.ends SAVM597

.subckt SAVM598 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2198 L=500e-9 W=3e-6
m2 net19 bl 0 0 N598 L=500e-9 W=3e-6
.ends SAVM598

.subckt SAVM599 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2199 L=500e-9 W=3e-6
m2 net19 bl 0 0 N599 L=500e-9 W=3e-6
.ends SAVM599

.subckt SAVM600 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2200 L=500e-9 W=3e-6
m2 net19 bl 0 0 N600 L=500e-9 W=3e-6
.ends SAVM600

.subckt SAVM601 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2201 L=500e-9 W=3e-6
m2 net19 bl 0 0 N601 L=500e-9 W=3e-6
.ends SAVM601

.subckt SAVM602 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2202 L=500e-9 W=3e-6
m2 net19 bl 0 0 N602 L=500e-9 W=3e-6
.ends SAVM602

.subckt SAVM603 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2203 L=500e-9 W=3e-6
m2 net19 bl 0 0 N603 L=500e-9 W=3e-6
.ends SAVM603

.subckt SAVM604 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2204 L=500e-9 W=3e-6
m2 net19 bl 0 0 N604 L=500e-9 W=3e-6
.ends SAVM604

.subckt SAVM605 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2205 L=500e-9 W=3e-6
m2 net19 bl 0 0 N605 L=500e-9 W=3e-6
.ends SAVM605

.subckt SAVM606 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2206 L=500e-9 W=3e-6
m2 net19 bl 0 0 N606 L=500e-9 W=3e-6
.ends SAVM606

.subckt SAVM607 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2207 L=500e-9 W=3e-6
m2 net19 bl 0 0 N607 L=500e-9 W=3e-6
.ends SAVM607

.subckt SAVM608 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2208 L=500e-9 W=3e-6
m2 net19 bl 0 0 N608 L=500e-9 W=3e-6
.ends SAVM608

.subckt SAVM609 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2209 L=500e-9 W=3e-6
m2 net19 bl 0 0 N609 L=500e-9 W=3e-6
.ends SAVM609

.subckt SAVM610 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2210 L=500e-9 W=3e-6
m2 net19 bl 0 0 N610 L=500e-9 W=3e-6
.ends SAVM610

.subckt SAVM611 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2211 L=500e-9 W=3e-6
m2 net19 bl 0 0 N611 L=500e-9 W=3e-6
.ends SAVM611

.subckt SAVM612 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2212 L=500e-9 W=3e-6
m2 net19 bl 0 0 N612 L=500e-9 W=3e-6
.ends SAVM612

.subckt SAVM613 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2213 L=500e-9 W=3e-6
m2 net19 bl 0 0 N613 L=500e-9 W=3e-6
.ends SAVM613

.subckt SAVM614 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2214 L=500e-9 W=3e-6
m2 net19 bl 0 0 N614 L=500e-9 W=3e-6
.ends SAVM614

.subckt SAVM615 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2215 L=500e-9 W=3e-6
m2 net19 bl 0 0 N615 L=500e-9 W=3e-6
.ends SAVM615

.subckt SAVM616 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2216 L=500e-9 W=3e-6
m2 net19 bl 0 0 N616 L=500e-9 W=3e-6
.ends SAVM616

.subckt SAVM617 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2217 L=500e-9 W=3e-6
m2 net19 bl 0 0 N617 L=500e-9 W=3e-6
.ends SAVM617

.subckt SAVM618 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2218 L=500e-9 W=3e-6
m2 net19 bl 0 0 N618 L=500e-9 W=3e-6
.ends SAVM618

.subckt SAVM619 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2219 L=500e-9 W=3e-6
m2 net19 bl 0 0 N619 L=500e-9 W=3e-6
.ends SAVM619

.subckt SAVM620 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2220 L=500e-9 W=3e-6
m2 net19 bl 0 0 N620 L=500e-9 W=3e-6
.ends SAVM620

.subckt SAVM621 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2221 L=500e-9 W=3e-6
m2 net19 bl 0 0 N621 L=500e-9 W=3e-6
.ends SAVM621

.subckt SAVM622 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2222 L=500e-9 W=3e-6
m2 net19 bl 0 0 N622 L=500e-9 W=3e-6
.ends SAVM622

.subckt SAVM623 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2223 L=500e-9 W=3e-6
m2 net19 bl 0 0 N623 L=500e-9 W=3e-6
.ends SAVM623

.subckt SAVM624 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2224 L=500e-9 W=3e-6
m2 net19 bl 0 0 N624 L=500e-9 W=3e-6
.ends SAVM624

.subckt SAVM625 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2225 L=500e-9 W=3e-6
m2 net19 bl 0 0 N625 L=500e-9 W=3e-6
.ends SAVM625

.subckt SAVM626 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2226 L=500e-9 W=3e-6
m2 net19 bl 0 0 N626 L=500e-9 W=3e-6
.ends SAVM626

.subckt SAVM627 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2227 L=500e-9 W=3e-6
m2 net19 bl 0 0 N627 L=500e-9 W=3e-6
.ends SAVM627

.subckt SAVM628 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2228 L=500e-9 W=3e-6
m2 net19 bl 0 0 N628 L=500e-9 W=3e-6
.ends SAVM628

.subckt SAVM629 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2229 L=500e-9 W=3e-6
m2 net19 bl 0 0 N629 L=500e-9 W=3e-6
.ends SAVM629

.subckt SAVM630 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2230 L=500e-9 W=3e-6
m2 net19 bl 0 0 N630 L=500e-9 W=3e-6
.ends SAVM630

.subckt SAVM631 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2231 L=500e-9 W=3e-6
m2 net19 bl 0 0 N631 L=500e-9 W=3e-6
.ends SAVM631

.subckt SAVM632 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2232 L=500e-9 W=3e-6
m2 net19 bl 0 0 N632 L=500e-9 W=3e-6
.ends SAVM632

.subckt SAVM633 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2233 L=500e-9 W=3e-6
m2 net19 bl 0 0 N633 L=500e-9 W=3e-6
.ends SAVM633

.subckt SAVM634 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2234 L=500e-9 W=3e-6
m2 net19 bl 0 0 N634 L=500e-9 W=3e-6
.ends SAVM634

.subckt SAVM635 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2235 L=500e-9 W=3e-6
m2 net19 bl 0 0 N635 L=500e-9 W=3e-6
.ends SAVM635

.subckt SAVM636 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2236 L=500e-9 W=3e-6
m2 net19 bl 0 0 N636 L=500e-9 W=3e-6
.ends SAVM636

.subckt SAVM637 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2237 L=500e-9 W=3e-6
m2 net19 bl 0 0 N637 L=500e-9 W=3e-6
.ends SAVM637

.subckt SAVM638 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2238 L=500e-9 W=3e-6
m2 net19 bl 0 0 N638 L=500e-9 W=3e-6
.ends SAVM638

.subckt SAVM639 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2239 L=500e-9 W=3e-6
m2 net19 bl 0 0 N639 L=500e-9 W=3e-6
.ends SAVM639

.subckt SAVM640 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2240 L=500e-9 W=3e-6
m2 net19 bl 0 0 N640 L=500e-9 W=3e-6
.ends SAVM640

.subckt SAVM641 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2241 L=500e-9 W=3e-6
m2 net19 bl 0 0 N641 L=500e-9 W=3e-6
.ends SAVM641

.subckt SAVM642 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2242 L=500e-9 W=3e-6
m2 net19 bl 0 0 N642 L=500e-9 W=3e-6
.ends SAVM642

.subckt SAVM643 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2243 L=500e-9 W=3e-6
m2 net19 bl 0 0 N643 L=500e-9 W=3e-6
.ends SAVM643

.subckt SAVM644 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2244 L=500e-9 W=3e-6
m2 net19 bl 0 0 N644 L=500e-9 W=3e-6
.ends SAVM644

.subckt SAVM645 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2245 L=500e-9 W=3e-6
m2 net19 bl 0 0 N645 L=500e-9 W=3e-6
.ends SAVM645

.subckt SAVM646 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2246 L=500e-9 W=3e-6
m2 net19 bl 0 0 N646 L=500e-9 W=3e-6
.ends SAVM646

.subckt SAVM647 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2247 L=500e-9 W=3e-6
m2 net19 bl 0 0 N647 L=500e-9 W=3e-6
.ends SAVM647

.subckt SAVM648 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2248 L=500e-9 W=3e-6
m2 net19 bl 0 0 N648 L=500e-9 W=3e-6
.ends SAVM648

.subckt SAVM649 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2249 L=500e-9 W=3e-6
m2 net19 bl 0 0 N649 L=500e-9 W=3e-6
.ends SAVM649

.subckt SAVM650 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2250 L=500e-9 W=3e-6
m2 net19 bl 0 0 N650 L=500e-9 W=3e-6
.ends SAVM650

.subckt SAVM651 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2251 L=500e-9 W=3e-6
m2 net19 bl 0 0 N651 L=500e-9 W=3e-6
.ends SAVM651

.subckt SAVM652 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2252 L=500e-9 W=3e-6
m2 net19 bl 0 0 N652 L=500e-9 W=3e-6
.ends SAVM652

.subckt SAVM653 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2253 L=500e-9 W=3e-6
m2 net19 bl 0 0 N653 L=500e-9 W=3e-6
.ends SAVM653

.subckt SAVM654 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2254 L=500e-9 W=3e-6
m2 net19 bl 0 0 N654 L=500e-9 W=3e-6
.ends SAVM654

.subckt SAVM655 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2255 L=500e-9 W=3e-6
m2 net19 bl 0 0 N655 L=500e-9 W=3e-6
.ends SAVM655

.subckt SAVM656 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2256 L=500e-9 W=3e-6
m2 net19 bl 0 0 N656 L=500e-9 W=3e-6
.ends SAVM656

.subckt SAVM657 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2257 L=500e-9 W=3e-6
m2 net19 bl 0 0 N657 L=500e-9 W=3e-6
.ends SAVM657

.subckt SAVM658 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2258 L=500e-9 W=3e-6
m2 net19 bl 0 0 N658 L=500e-9 W=3e-6
.ends SAVM658

.subckt SAVM659 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2259 L=500e-9 W=3e-6
m2 net19 bl 0 0 N659 L=500e-9 W=3e-6
.ends SAVM659

.subckt SAVM660 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2260 L=500e-9 W=3e-6
m2 net19 bl 0 0 N660 L=500e-9 W=3e-6
.ends SAVM660

.subckt SAVM661 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2261 L=500e-9 W=3e-6
m2 net19 bl 0 0 N661 L=500e-9 W=3e-6
.ends SAVM661

.subckt SAVM662 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2262 L=500e-9 W=3e-6
m2 net19 bl 0 0 N662 L=500e-9 W=3e-6
.ends SAVM662

.subckt SAVM663 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2263 L=500e-9 W=3e-6
m2 net19 bl 0 0 N663 L=500e-9 W=3e-6
.ends SAVM663

.subckt SAVM664 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2264 L=500e-9 W=3e-6
m2 net19 bl 0 0 N664 L=500e-9 W=3e-6
.ends SAVM664

.subckt SAVM665 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2265 L=500e-9 W=3e-6
m2 net19 bl 0 0 N665 L=500e-9 W=3e-6
.ends SAVM665

.subckt SAVM666 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2266 L=500e-9 W=3e-6
m2 net19 bl 0 0 N666 L=500e-9 W=3e-6
.ends SAVM666

.subckt SAVM667 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2267 L=500e-9 W=3e-6
m2 net19 bl 0 0 N667 L=500e-9 W=3e-6
.ends SAVM667

.subckt SAVM668 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2268 L=500e-9 W=3e-6
m2 net19 bl 0 0 N668 L=500e-9 W=3e-6
.ends SAVM668

.subckt SAVM669 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2269 L=500e-9 W=3e-6
m2 net19 bl 0 0 N669 L=500e-9 W=3e-6
.ends SAVM669

.subckt SAVM670 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2270 L=500e-9 W=3e-6
m2 net19 bl 0 0 N670 L=500e-9 W=3e-6
.ends SAVM670

.subckt SAVM671 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2271 L=500e-9 W=3e-6
m2 net19 bl 0 0 N671 L=500e-9 W=3e-6
.ends SAVM671

.subckt SAVM672 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2272 L=500e-9 W=3e-6
m2 net19 bl 0 0 N672 L=500e-9 W=3e-6
.ends SAVM672

.subckt SAVM673 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2273 L=500e-9 W=3e-6
m2 net19 bl 0 0 N673 L=500e-9 W=3e-6
.ends SAVM673

.subckt SAVM674 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2274 L=500e-9 W=3e-6
m2 net19 bl 0 0 N674 L=500e-9 W=3e-6
.ends SAVM674

.subckt SAVM675 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2275 L=500e-9 W=3e-6
m2 net19 bl 0 0 N675 L=500e-9 W=3e-6
.ends SAVM675

.subckt SAVM676 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2276 L=500e-9 W=3e-6
m2 net19 bl 0 0 N676 L=500e-9 W=3e-6
.ends SAVM676

.subckt SAVM677 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2277 L=500e-9 W=3e-6
m2 net19 bl 0 0 N677 L=500e-9 W=3e-6
.ends SAVM677

.subckt SAVM678 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2278 L=500e-9 W=3e-6
m2 net19 bl 0 0 N678 L=500e-9 W=3e-6
.ends SAVM678

.subckt SAVM679 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2279 L=500e-9 W=3e-6
m2 net19 bl 0 0 N679 L=500e-9 W=3e-6
.ends SAVM679

.subckt SAVM680 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2280 L=500e-9 W=3e-6
m2 net19 bl 0 0 N680 L=500e-9 W=3e-6
.ends SAVM680

.subckt SAVM681 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2281 L=500e-9 W=3e-6
m2 net19 bl 0 0 N681 L=500e-9 W=3e-6
.ends SAVM681

.subckt SAVM682 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2282 L=500e-9 W=3e-6
m2 net19 bl 0 0 N682 L=500e-9 W=3e-6
.ends SAVM682

.subckt SAVM683 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2283 L=500e-9 W=3e-6
m2 net19 bl 0 0 N683 L=500e-9 W=3e-6
.ends SAVM683

.subckt SAVM684 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2284 L=500e-9 W=3e-6
m2 net19 bl 0 0 N684 L=500e-9 W=3e-6
.ends SAVM684

.subckt SAVM685 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2285 L=500e-9 W=3e-6
m2 net19 bl 0 0 N685 L=500e-9 W=3e-6
.ends SAVM685

.subckt SAVM686 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2286 L=500e-9 W=3e-6
m2 net19 bl 0 0 N686 L=500e-9 W=3e-6
.ends SAVM686

.subckt SAVM687 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2287 L=500e-9 W=3e-6
m2 net19 bl 0 0 N687 L=500e-9 W=3e-6
.ends SAVM687

.subckt SAVM688 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2288 L=500e-9 W=3e-6
m2 net19 bl 0 0 N688 L=500e-9 W=3e-6
.ends SAVM688

.subckt SAVM689 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2289 L=500e-9 W=3e-6
m2 net19 bl 0 0 N689 L=500e-9 W=3e-6
.ends SAVM689

.subckt SAVM690 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2290 L=500e-9 W=3e-6
m2 net19 bl 0 0 N690 L=500e-9 W=3e-6
.ends SAVM690

.subckt SAVM691 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2291 L=500e-9 W=3e-6
m2 net19 bl 0 0 N691 L=500e-9 W=3e-6
.ends SAVM691

.subckt SAVM692 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2292 L=500e-9 W=3e-6
m2 net19 bl 0 0 N692 L=500e-9 W=3e-6
.ends SAVM692

.subckt SAVM693 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2293 L=500e-9 W=3e-6
m2 net19 bl 0 0 N693 L=500e-9 W=3e-6
.ends SAVM693

.subckt SAVM694 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2294 L=500e-9 W=3e-6
m2 net19 bl 0 0 N694 L=500e-9 W=3e-6
.ends SAVM694

.subckt SAVM695 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2295 L=500e-9 W=3e-6
m2 net19 bl 0 0 N695 L=500e-9 W=3e-6
.ends SAVM695

.subckt SAVM696 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2296 L=500e-9 W=3e-6
m2 net19 bl 0 0 N696 L=500e-9 W=3e-6
.ends SAVM696

.subckt SAVM697 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2297 L=500e-9 W=3e-6
m2 net19 bl 0 0 N697 L=500e-9 W=3e-6
.ends SAVM697

.subckt SAVM698 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2298 L=500e-9 W=3e-6
m2 net19 bl 0 0 N698 L=500e-9 W=3e-6
.ends SAVM698

.subckt SAVM699 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2299 L=500e-9 W=3e-6
m2 net19 bl 0 0 N699 L=500e-9 W=3e-6
.ends SAVM699

.subckt SAVM700 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2300 L=500e-9 W=3e-6
m2 net19 bl 0 0 N700 L=500e-9 W=3e-6
.ends SAVM700

.subckt SAVM701 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2301 L=500e-9 W=3e-6
m2 net19 bl 0 0 N701 L=500e-9 W=3e-6
.ends SAVM701

.subckt SAVM702 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2302 L=500e-9 W=3e-6
m2 net19 bl 0 0 N702 L=500e-9 W=3e-6
.ends SAVM702

.subckt SAVM703 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2303 L=500e-9 W=3e-6
m2 net19 bl 0 0 N703 L=500e-9 W=3e-6
.ends SAVM703

.subckt SAVM704 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2304 L=500e-9 W=3e-6
m2 net19 bl 0 0 N704 L=500e-9 W=3e-6
.ends SAVM704

.subckt SAVM705 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2305 L=500e-9 W=3e-6
m2 net19 bl 0 0 N705 L=500e-9 W=3e-6
.ends SAVM705

.subckt SAVM706 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2306 L=500e-9 W=3e-6
m2 net19 bl 0 0 N706 L=500e-9 W=3e-6
.ends SAVM706

.subckt SAVM707 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2307 L=500e-9 W=3e-6
m2 net19 bl 0 0 N707 L=500e-9 W=3e-6
.ends SAVM707

.subckt SAVM708 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2308 L=500e-9 W=3e-6
m2 net19 bl 0 0 N708 L=500e-9 W=3e-6
.ends SAVM708

.subckt SAVM709 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2309 L=500e-9 W=3e-6
m2 net19 bl 0 0 N709 L=500e-9 W=3e-6
.ends SAVM709

.subckt SAVM710 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2310 L=500e-9 W=3e-6
m2 net19 bl 0 0 N710 L=500e-9 W=3e-6
.ends SAVM710

.subckt SAVM711 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2311 L=500e-9 W=3e-6
m2 net19 bl 0 0 N711 L=500e-9 W=3e-6
.ends SAVM711

.subckt SAVM712 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2312 L=500e-9 W=3e-6
m2 net19 bl 0 0 N712 L=500e-9 W=3e-6
.ends SAVM712

.subckt SAVM713 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2313 L=500e-9 W=3e-6
m2 net19 bl 0 0 N713 L=500e-9 W=3e-6
.ends SAVM713

.subckt SAVM714 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2314 L=500e-9 W=3e-6
m2 net19 bl 0 0 N714 L=500e-9 W=3e-6
.ends SAVM714

.subckt SAVM715 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2315 L=500e-9 W=3e-6
m2 net19 bl 0 0 N715 L=500e-9 W=3e-6
.ends SAVM715

.subckt SAVM716 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2316 L=500e-9 W=3e-6
m2 net19 bl 0 0 N716 L=500e-9 W=3e-6
.ends SAVM716

.subckt SAVM717 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2317 L=500e-9 W=3e-6
m2 net19 bl 0 0 N717 L=500e-9 W=3e-6
.ends SAVM717

.subckt SAVM718 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2318 L=500e-9 W=3e-6
m2 net19 bl 0 0 N718 L=500e-9 W=3e-6
.ends SAVM718

.subckt SAVM719 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2319 L=500e-9 W=3e-6
m2 net19 bl 0 0 N719 L=500e-9 W=3e-6
.ends SAVM719

.subckt SAVM720 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2320 L=500e-9 W=3e-6
m2 net19 bl 0 0 N720 L=500e-9 W=3e-6
.ends SAVM720

.subckt SAVM721 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2321 L=500e-9 W=3e-6
m2 net19 bl 0 0 N721 L=500e-9 W=3e-6
.ends SAVM721

.subckt SAVM722 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2322 L=500e-9 W=3e-6
m2 net19 bl 0 0 N722 L=500e-9 W=3e-6
.ends SAVM722

.subckt SAVM723 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2323 L=500e-9 W=3e-6
m2 net19 bl 0 0 N723 L=500e-9 W=3e-6
.ends SAVM723

.subckt SAVM724 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2324 L=500e-9 W=3e-6
m2 net19 bl 0 0 N724 L=500e-9 W=3e-6
.ends SAVM724

.subckt SAVM725 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2325 L=500e-9 W=3e-6
m2 net19 bl 0 0 N725 L=500e-9 W=3e-6
.ends SAVM725

.subckt SAVM726 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2326 L=500e-9 W=3e-6
m2 net19 bl 0 0 N726 L=500e-9 W=3e-6
.ends SAVM726

.subckt SAVM727 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2327 L=500e-9 W=3e-6
m2 net19 bl 0 0 N727 L=500e-9 W=3e-6
.ends SAVM727

.subckt SAVM728 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2328 L=500e-9 W=3e-6
m2 net19 bl 0 0 N728 L=500e-9 W=3e-6
.ends SAVM728

.subckt SAVM729 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2329 L=500e-9 W=3e-6
m2 net19 bl 0 0 N729 L=500e-9 W=3e-6
.ends SAVM729

.subckt SAVM730 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2330 L=500e-9 W=3e-6
m2 net19 bl 0 0 N730 L=500e-9 W=3e-6
.ends SAVM730

.subckt SAVM731 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2331 L=500e-9 W=3e-6
m2 net19 bl 0 0 N731 L=500e-9 W=3e-6
.ends SAVM731

.subckt SAVM732 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2332 L=500e-9 W=3e-6
m2 net19 bl 0 0 N732 L=500e-9 W=3e-6
.ends SAVM732

.subckt SAVM733 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2333 L=500e-9 W=3e-6
m2 net19 bl 0 0 N733 L=500e-9 W=3e-6
.ends SAVM733

.subckt SAVM734 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2334 L=500e-9 W=3e-6
m2 net19 bl 0 0 N734 L=500e-9 W=3e-6
.ends SAVM734

.subckt SAVM735 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2335 L=500e-9 W=3e-6
m2 net19 bl 0 0 N735 L=500e-9 W=3e-6
.ends SAVM735

.subckt SAVM736 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2336 L=500e-9 W=3e-6
m2 net19 bl 0 0 N736 L=500e-9 W=3e-6
.ends SAVM736

.subckt SAVM737 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2337 L=500e-9 W=3e-6
m2 net19 bl 0 0 N737 L=500e-9 W=3e-6
.ends SAVM737

.subckt SAVM738 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2338 L=500e-9 W=3e-6
m2 net19 bl 0 0 N738 L=500e-9 W=3e-6
.ends SAVM738

.subckt SAVM739 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2339 L=500e-9 W=3e-6
m2 net19 bl 0 0 N739 L=500e-9 W=3e-6
.ends SAVM739

.subckt SAVM740 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2340 L=500e-9 W=3e-6
m2 net19 bl 0 0 N740 L=500e-9 W=3e-6
.ends SAVM740

.subckt SAVM741 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2341 L=500e-9 W=3e-6
m2 net19 bl 0 0 N741 L=500e-9 W=3e-6
.ends SAVM741

.subckt SAVM742 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2342 L=500e-9 W=3e-6
m2 net19 bl 0 0 N742 L=500e-9 W=3e-6
.ends SAVM742

.subckt SAVM743 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2343 L=500e-9 W=3e-6
m2 net19 bl 0 0 N743 L=500e-9 W=3e-6
.ends SAVM743

.subckt SAVM744 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2344 L=500e-9 W=3e-6
m2 net19 bl 0 0 N744 L=500e-9 W=3e-6
.ends SAVM744

.subckt SAVM745 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2345 L=500e-9 W=3e-6
m2 net19 bl 0 0 N745 L=500e-9 W=3e-6
.ends SAVM745

.subckt SAVM746 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2346 L=500e-9 W=3e-6
m2 net19 bl 0 0 N746 L=500e-9 W=3e-6
.ends SAVM746

.subckt SAVM747 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2347 L=500e-9 W=3e-6
m2 net19 bl 0 0 N747 L=500e-9 W=3e-6
.ends SAVM747

.subckt SAVM748 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2348 L=500e-9 W=3e-6
m2 net19 bl 0 0 N748 L=500e-9 W=3e-6
.ends SAVM748

.subckt SAVM749 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2349 L=500e-9 W=3e-6
m2 net19 bl 0 0 N749 L=500e-9 W=3e-6
.ends SAVM749

.subckt SAVM750 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2350 L=500e-9 W=3e-6
m2 net19 bl 0 0 N750 L=500e-9 W=3e-6
.ends SAVM750

.subckt SAVM751 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2351 L=500e-9 W=3e-6
m2 net19 bl 0 0 N751 L=500e-9 W=3e-6
.ends SAVM751

.subckt SAVM752 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2352 L=500e-9 W=3e-6
m2 net19 bl 0 0 N752 L=500e-9 W=3e-6
.ends SAVM752

.subckt SAVM753 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2353 L=500e-9 W=3e-6
m2 net19 bl 0 0 N753 L=500e-9 W=3e-6
.ends SAVM753

.subckt SAVM754 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2354 L=500e-9 W=3e-6
m2 net19 bl 0 0 N754 L=500e-9 W=3e-6
.ends SAVM754

.subckt SAVM755 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2355 L=500e-9 W=3e-6
m2 net19 bl 0 0 N755 L=500e-9 W=3e-6
.ends SAVM755

.subckt SAVM756 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2356 L=500e-9 W=3e-6
m2 net19 bl 0 0 N756 L=500e-9 W=3e-6
.ends SAVM756

.subckt SAVM757 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2357 L=500e-9 W=3e-6
m2 net19 bl 0 0 N757 L=500e-9 W=3e-6
.ends SAVM757

.subckt SAVM758 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2358 L=500e-9 W=3e-6
m2 net19 bl 0 0 N758 L=500e-9 W=3e-6
.ends SAVM758

.subckt SAVM759 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2359 L=500e-9 W=3e-6
m2 net19 bl 0 0 N759 L=500e-9 W=3e-6
.ends SAVM759

.subckt SAVM760 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2360 L=500e-9 W=3e-6
m2 net19 bl 0 0 N760 L=500e-9 W=3e-6
.ends SAVM760

.subckt SAVM761 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2361 L=500e-9 W=3e-6
m2 net19 bl 0 0 N761 L=500e-9 W=3e-6
.ends SAVM761

.subckt SAVM762 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2362 L=500e-9 W=3e-6
m2 net19 bl 0 0 N762 L=500e-9 W=3e-6
.ends SAVM762

.subckt SAVM763 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2363 L=500e-9 W=3e-6
m2 net19 bl 0 0 N763 L=500e-9 W=3e-6
.ends SAVM763

.subckt SAVM764 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2364 L=500e-9 W=3e-6
m2 net19 bl 0 0 N764 L=500e-9 W=3e-6
.ends SAVM764

.subckt SAVM765 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2365 L=500e-9 W=3e-6
m2 net19 bl 0 0 N765 L=500e-9 W=3e-6
.ends SAVM765

.subckt SAVM766 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2366 L=500e-9 W=3e-6
m2 net19 bl 0 0 N766 L=500e-9 W=3e-6
.ends SAVM766

.subckt SAVM767 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2367 L=500e-9 W=3e-6
m2 net19 bl 0 0 N767 L=500e-9 W=3e-6
.ends SAVM767

.subckt SAVM768 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2368 L=500e-9 W=3e-6
m2 net19 bl 0 0 N768 L=500e-9 W=3e-6
.ends SAVM768

.subckt SAVM769 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2369 L=500e-9 W=3e-6
m2 net19 bl 0 0 N769 L=500e-9 W=3e-6
.ends SAVM769

.subckt SAVM770 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2370 L=500e-9 W=3e-6
m2 net19 bl 0 0 N770 L=500e-9 W=3e-6
.ends SAVM770

.subckt SAVM771 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2371 L=500e-9 W=3e-6
m2 net19 bl 0 0 N771 L=500e-9 W=3e-6
.ends SAVM771

.subckt SAVM772 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2372 L=500e-9 W=3e-6
m2 net19 bl 0 0 N772 L=500e-9 W=3e-6
.ends SAVM772

.subckt SAVM773 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2373 L=500e-9 W=3e-6
m2 net19 bl 0 0 N773 L=500e-9 W=3e-6
.ends SAVM773

.subckt SAVM774 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2374 L=500e-9 W=3e-6
m2 net19 bl 0 0 N774 L=500e-9 W=3e-6
.ends SAVM774

.subckt SAVM775 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2375 L=500e-9 W=3e-6
m2 net19 bl 0 0 N775 L=500e-9 W=3e-6
.ends SAVM775

.subckt SAVM776 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2376 L=500e-9 W=3e-6
m2 net19 bl 0 0 N776 L=500e-9 W=3e-6
.ends SAVM776

.subckt SAVM777 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2377 L=500e-9 W=3e-6
m2 net19 bl 0 0 N777 L=500e-9 W=3e-6
.ends SAVM777

.subckt SAVM778 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2378 L=500e-9 W=3e-6
m2 net19 bl 0 0 N778 L=500e-9 W=3e-6
.ends SAVM778

.subckt SAVM779 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2379 L=500e-9 W=3e-6
m2 net19 bl 0 0 N779 L=500e-9 W=3e-6
.ends SAVM779

.subckt SAVM780 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2380 L=500e-9 W=3e-6
m2 net19 bl 0 0 N780 L=500e-9 W=3e-6
.ends SAVM780

.subckt SAVM781 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2381 L=500e-9 W=3e-6
m2 net19 bl 0 0 N781 L=500e-9 W=3e-6
.ends SAVM781

.subckt SAVM782 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2382 L=500e-9 W=3e-6
m2 net19 bl 0 0 N782 L=500e-9 W=3e-6
.ends SAVM782

.subckt SAVM783 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2383 L=500e-9 W=3e-6
m2 net19 bl 0 0 N783 L=500e-9 W=3e-6
.ends SAVM783

.subckt SAVM784 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2384 L=500e-9 W=3e-6
m2 net19 bl 0 0 N784 L=500e-9 W=3e-6
.ends SAVM784

.subckt SAVM785 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2385 L=500e-9 W=3e-6
m2 net19 bl 0 0 N785 L=500e-9 W=3e-6
.ends SAVM785

.subckt SAVM786 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2386 L=500e-9 W=3e-6
m2 net19 bl 0 0 N786 L=500e-9 W=3e-6
.ends SAVM786

.subckt SAVM787 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2387 L=500e-9 W=3e-6
m2 net19 bl 0 0 N787 L=500e-9 W=3e-6
.ends SAVM787

.subckt SAVM788 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2388 L=500e-9 W=3e-6
m2 net19 bl 0 0 N788 L=500e-9 W=3e-6
.ends SAVM788

.subckt SAVM789 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2389 L=500e-9 W=3e-6
m2 net19 bl 0 0 N789 L=500e-9 W=3e-6
.ends SAVM789

.subckt SAVM790 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2390 L=500e-9 W=3e-6
m2 net19 bl 0 0 N790 L=500e-9 W=3e-6
.ends SAVM790

.subckt SAVM791 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2391 L=500e-9 W=3e-6
m2 net19 bl 0 0 N791 L=500e-9 W=3e-6
.ends SAVM791

.subckt SAVM792 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2392 L=500e-9 W=3e-6
m2 net19 bl 0 0 N792 L=500e-9 W=3e-6
.ends SAVM792

.subckt SAVM793 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2393 L=500e-9 W=3e-6
m2 net19 bl 0 0 N793 L=500e-9 W=3e-6
.ends SAVM793

.subckt SAVM794 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2394 L=500e-9 W=3e-6
m2 net19 bl 0 0 N794 L=500e-9 W=3e-6
.ends SAVM794

.subckt SAVM795 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2395 L=500e-9 W=3e-6
m2 net19 bl 0 0 N795 L=500e-9 W=3e-6
.ends SAVM795

.subckt SAVM796 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2396 L=500e-9 W=3e-6
m2 net19 bl 0 0 N796 L=500e-9 W=3e-6
.ends SAVM796

.subckt SAVM797 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2397 L=500e-9 W=3e-6
m2 net19 bl 0 0 N797 L=500e-9 W=3e-6
.ends SAVM797

.subckt SAVM798 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2398 L=500e-9 W=3e-6
m2 net19 bl 0 0 N798 L=500e-9 W=3e-6
.ends SAVM798

.subckt SAVM799 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2399 L=500e-9 W=3e-6
m2 net19 bl 0 0 N799 L=500e-9 W=3e-6
.ends SAVM799

.subckt SAVM800 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2400 L=500e-9 W=3e-6
m2 net19 bl 0 0 N800 L=500e-9 W=3e-6
.ends SAVM800

.subckt SAVM801 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2401 L=500e-9 W=3e-6
m2 net19 bl 0 0 N801 L=500e-9 W=3e-6
.ends SAVM801

.subckt SAVM802 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2402 L=500e-9 W=3e-6
m2 net19 bl 0 0 N802 L=500e-9 W=3e-6
.ends SAVM802

.subckt SAVM803 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2403 L=500e-9 W=3e-6
m2 net19 bl 0 0 N803 L=500e-9 W=3e-6
.ends SAVM803

.subckt SAVM804 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2404 L=500e-9 W=3e-6
m2 net19 bl 0 0 N804 L=500e-9 W=3e-6
.ends SAVM804

.subckt SAVM805 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2405 L=500e-9 W=3e-6
m2 net19 bl 0 0 N805 L=500e-9 W=3e-6
.ends SAVM805

.subckt SAVM806 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2406 L=500e-9 W=3e-6
m2 net19 bl 0 0 N806 L=500e-9 W=3e-6
.ends SAVM806

.subckt SAVM807 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2407 L=500e-9 W=3e-6
m2 net19 bl 0 0 N807 L=500e-9 W=3e-6
.ends SAVM807

.subckt SAVM808 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2408 L=500e-9 W=3e-6
m2 net19 bl 0 0 N808 L=500e-9 W=3e-6
.ends SAVM808

.subckt SAVM809 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2409 L=500e-9 W=3e-6
m2 net19 bl 0 0 N809 L=500e-9 W=3e-6
.ends SAVM809

.subckt SAVM810 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2410 L=500e-9 W=3e-6
m2 net19 bl 0 0 N810 L=500e-9 W=3e-6
.ends SAVM810

.subckt SAVM811 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2411 L=500e-9 W=3e-6
m2 net19 bl 0 0 N811 L=500e-9 W=3e-6
.ends SAVM811

.subckt SAVM812 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2412 L=500e-9 W=3e-6
m2 net19 bl 0 0 N812 L=500e-9 W=3e-6
.ends SAVM812

.subckt SAVM813 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2413 L=500e-9 W=3e-6
m2 net19 bl 0 0 N813 L=500e-9 W=3e-6
.ends SAVM813

.subckt SAVM814 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2414 L=500e-9 W=3e-6
m2 net19 bl 0 0 N814 L=500e-9 W=3e-6
.ends SAVM814

.subckt SAVM815 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2415 L=500e-9 W=3e-6
m2 net19 bl 0 0 N815 L=500e-9 W=3e-6
.ends SAVM815

.subckt SAVM816 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2416 L=500e-9 W=3e-6
m2 net19 bl 0 0 N816 L=500e-9 W=3e-6
.ends SAVM816

.subckt SAVM817 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2417 L=500e-9 W=3e-6
m2 net19 bl 0 0 N817 L=500e-9 W=3e-6
.ends SAVM817

.subckt SAVM818 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2418 L=500e-9 W=3e-6
m2 net19 bl 0 0 N818 L=500e-9 W=3e-6
.ends SAVM818

.subckt SAVM819 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2419 L=500e-9 W=3e-6
m2 net19 bl 0 0 N819 L=500e-9 W=3e-6
.ends SAVM819

.subckt SAVM820 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2420 L=500e-9 W=3e-6
m2 net19 bl 0 0 N820 L=500e-9 W=3e-6
.ends SAVM820

.subckt SAVM821 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2421 L=500e-9 W=3e-6
m2 net19 bl 0 0 N821 L=500e-9 W=3e-6
.ends SAVM821

.subckt SAVM822 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2422 L=500e-9 W=3e-6
m2 net19 bl 0 0 N822 L=500e-9 W=3e-6
.ends SAVM822

.subckt SAVM823 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2423 L=500e-9 W=3e-6
m2 net19 bl 0 0 N823 L=500e-9 W=3e-6
.ends SAVM823

.subckt SAVM824 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2424 L=500e-9 W=3e-6
m2 net19 bl 0 0 N824 L=500e-9 W=3e-6
.ends SAVM824

.subckt SAVM825 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2425 L=500e-9 W=3e-6
m2 net19 bl 0 0 N825 L=500e-9 W=3e-6
.ends SAVM825

.subckt SAVM826 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2426 L=500e-9 W=3e-6
m2 net19 bl 0 0 N826 L=500e-9 W=3e-6
.ends SAVM826

.subckt SAVM827 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2427 L=500e-9 W=3e-6
m2 net19 bl 0 0 N827 L=500e-9 W=3e-6
.ends SAVM827

.subckt SAVM828 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2428 L=500e-9 W=3e-6
m2 net19 bl 0 0 N828 L=500e-9 W=3e-6
.ends SAVM828

.subckt SAVM829 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2429 L=500e-9 W=3e-6
m2 net19 bl 0 0 N829 L=500e-9 W=3e-6
.ends SAVM829

.subckt SAVM830 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2430 L=500e-9 W=3e-6
m2 net19 bl 0 0 N830 L=500e-9 W=3e-6
.ends SAVM830

.subckt SAVM831 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2431 L=500e-9 W=3e-6
m2 net19 bl 0 0 N831 L=500e-9 W=3e-6
.ends SAVM831

.subckt SAVM832 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2432 L=500e-9 W=3e-6
m2 net19 bl 0 0 N832 L=500e-9 W=3e-6
.ends SAVM832

.subckt SAVM833 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2433 L=500e-9 W=3e-6
m2 net19 bl 0 0 N833 L=500e-9 W=3e-6
.ends SAVM833

.subckt SAVM834 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2434 L=500e-9 W=3e-6
m2 net19 bl 0 0 N834 L=500e-9 W=3e-6
.ends SAVM834

.subckt SAVM835 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2435 L=500e-9 W=3e-6
m2 net19 bl 0 0 N835 L=500e-9 W=3e-6
.ends SAVM835

.subckt SAVM836 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2436 L=500e-9 W=3e-6
m2 net19 bl 0 0 N836 L=500e-9 W=3e-6
.ends SAVM836

.subckt SAVM837 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2437 L=500e-9 W=3e-6
m2 net19 bl 0 0 N837 L=500e-9 W=3e-6
.ends SAVM837

.subckt SAVM838 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2438 L=500e-9 W=3e-6
m2 net19 bl 0 0 N838 L=500e-9 W=3e-6
.ends SAVM838

.subckt SAVM839 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2439 L=500e-9 W=3e-6
m2 net19 bl 0 0 N839 L=500e-9 W=3e-6
.ends SAVM839

.subckt SAVM840 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2440 L=500e-9 W=3e-6
m2 net19 bl 0 0 N840 L=500e-9 W=3e-6
.ends SAVM840

.subckt SAVM841 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2441 L=500e-9 W=3e-6
m2 net19 bl 0 0 N841 L=500e-9 W=3e-6
.ends SAVM841

.subckt SAVM842 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2442 L=500e-9 W=3e-6
m2 net19 bl 0 0 N842 L=500e-9 W=3e-6
.ends SAVM842

.subckt SAVM843 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2443 L=500e-9 W=3e-6
m2 net19 bl 0 0 N843 L=500e-9 W=3e-6
.ends SAVM843

.subckt SAVM844 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2444 L=500e-9 W=3e-6
m2 net19 bl 0 0 N844 L=500e-9 W=3e-6
.ends SAVM844

.subckt SAVM845 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2445 L=500e-9 W=3e-6
m2 net19 bl 0 0 N845 L=500e-9 W=3e-6
.ends SAVM845

.subckt SAVM846 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2446 L=500e-9 W=3e-6
m2 net19 bl 0 0 N846 L=500e-9 W=3e-6
.ends SAVM846

.subckt SAVM847 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2447 L=500e-9 W=3e-6
m2 net19 bl 0 0 N847 L=500e-9 W=3e-6
.ends SAVM847

.subckt SAVM848 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2448 L=500e-9 W=3e-6
m2 net19 bl 0 0 N848 L=500e-9 W=3e-6
.ends SAVM848

.subckt SAVM849 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2449 L=500e-9 W=3e-6
m2 net19 bl 0 0 N849 L=500e-9 W=3e-6
.ends SAVM849

.subckt SAVM850 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2450 L=500e-9 W=3e-6
m2 net19 bl 0 0 N850 L=500e-9 W=3e-6
.ends SAVM850

.subckt SAVM851 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2451 L=500e-9 W=3e-6
m2 net19 bl 0 0 N851 L=500e-9 W=3e-6
.ends SAVM851

.subckt SAVM852 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2452 L=500e-9 W=3e-6
m2 net19 bl 0 0 N852 L=500e-9 W=3e-6
.ends SAVM852

.subckt SAVM853 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2453 L=500e-9 W=3e-6
m2 net19 bl 0 0 N853 L=500e-9 W=3e-6
.ends SAVM853

.subckt SAVM854 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2454 L=500e-9 W=3e-6
m2 net19 bl 0 0 N854 L=500e-9 W=3e-6
.ends SAVM854

.subckt SAVM855 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2455 L=500e-9 W=3e-6
m2 net19 bl 0 0 N855 L=500e-9 W=3e-6
.ends SAVM855

.subckt SAVM856 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2456 L=500e-9 W=3e-6
m2 net19 bl 0 0 N856 L=500e-9 W=3e-6
.ends SAVM856

.subckt SAVM857 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2457 L=500e-9 W=3e-6
m2 net19 bl 0 0 N857 L=500e-9 W=3e-6
.ends SAVM857

.subckt SAVM858 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2458 L=500e-9 W=3e-6
m2 net19 bl 0 0 N858 L=500e-9 W=3e-6
.ends SAVM858

.subckt SAVM859 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2459 L=500e-9 W=3e-6
m2 net19 bl 0 0 N859 L=500e-9 W=3e-6
.ends SAVM859

.subckt SAVM860 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2460 L=500e-9 W=3e-6
m2 net19 bl 0 0 N860 L=500e-9 W=3e-6
.ends SAVM860

.subckt SAVM861 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2461 L=500e-9 W=3e-6
m2 net19 bl 0 0 N861 L=500e-9 W=3e-6
.ends SAVM861

.subckt SAVM862 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2462 L=500e-9 W=3e-6
m2 net19 bl 0 0 N862 L=500e-9 W=3e-6
.ends SAVM862

.subckt SAVM863 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2463 L=500e-9 W=3e-6
m2 net19 bl 0 0 N863 L=500e-9 W=3e-6
.ends SAVM863

.subckt SAVM864 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2464 L=500e-9 W=3e-6
m2 net19 bl 0 0 N864 L=500e-9 W=3e-6
.ends SAVM864

.subckt SAVM865 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2465 L=500e-9 W=3e-6
m2 net19 bl 0 0 N865 L=500e-9 W=3e-6
.ends SAVM865

.subckt SAVM866 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2466 L=500e-9 W=3e-6
m2 net19 bl 0 0 N866 L=500e-9 W=3e-6
.ends SAVM866

.subckt SAVM867 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2467 L=500e-9 W=3e-6
m2 net19 bl 0 0 N867 L=500e-9 W=3e-6
.ends SAVM867

.subckt SAVM868 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2468 L=500e-9 W=3e-6
m2 net19 bl 0 0 N868 L=500e-9 W=3e-6
.ends SAVM868

.subckt SAVM869 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2469 L=500e-9 W=3e-6
m2 net19 bl 0 0 N869 L=500e-9 W=3e-6
.ends SAVM869

.subckt SAVM870 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2470 L=500e-9 W=3e-6
m2 net19 bl 0 0 N870 L=500e-9 W=3e-6
.ends SAVM870

.subckt SAVM871 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2471 L=500e-9 W=3e-6
m2 net19 bl 0 0 N871 L=500e-9 W=3e-6
.ends SAVM871

.subckt SAVM872 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2472 L=500e-9 W=3e-6
m2 net19 bl 0 0 N872 L=500e-9 W=3e-6
.ends SAVM872

.subckt SAVM873 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2473 L=500e-9 W=3e-6
m2 net19 bl 0 0 N873 L=500e-9 W=3e-6
.ends SAVM873

.subckt SAVM874 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2474 L=500e-9 W=3e-6
m2 net19 bl 0 0 N874 L=500e-9 W=3e-6
.ends SAVM874

.subckt SAVM875 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2475 L=500e-9 W=3e-6
m2 net19 bl 0 0 N875 L=500e-9 W=3e-6
.ends SAVM875

.subckt SAVM876 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2476 L=500e-9 W=3e-6
m2 net19 bl 0 0 N876 L=500e-9 W=3e-6
.ends SAVM876

.subckt SAVM877 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2477 L=500e-9 W=3e-6
m2 net19 bl 0 0 N877 L=500e-9 W=3e-6
.ends SAVM877

.subckt SAVM878 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2478 L=500e-9 W=3e-6
m2 net19 bl 0 0 N878 L=500e-9 W=3e-6
.ends SAVM878

.subckt SAVM879 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2479 L=500e-9 W=3e-6
m2 net19 bl 0 0 N879 L=500e-9 W=3e-6
.ends SAVM879

.subckt SAVM880 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2480 L=500e-9 W=3e-6
m2 net19 bl 0 0 N880 L=500e-9 W=3e-6
.ends SAVM880

.subckt SAVM881 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2481 L=500e-9 W=3e-6
m2 net19 bl 0 0 N881 L=500e-9 W=3e-6
.ends SAVM881

.subckt SAVM882 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2482 L=500e-9 W=3e-6
m2 net19 bl 0 0 N882 L=500e-9 W=3e-6
.ends SAVM882

.subckt SAVM883 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2483 L=500e-9 W=3e-6
m2 net19 bl 0 0 N883 L=500e-9 W=3e-6
.ends SAVM883

.subckt SAVM884 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2484 L=500e-9 W=3e-6
m2 net19 bl 0 0 N884 L=500e-9 W=3e-6
.ends SAVM884

.subckt SAVM885 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2485 L=500e-9 W=3e-6
m2 net19 bl 0 0 N885 L=500e-9 W=3e-6
.ends SAVM885

.subckt SAVM886 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2486 L=500e-9 W=3e-6
m2 net19 bl 0 0 N886 L=500e-9 W=3e-6
.ends SAVM886

.subckt SAVM887 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2487 L=500e-9 W=3e-6
m2 net19 bl 0 0 N887 L=500e-9 W=3e-6
.ends SAVM887

.subckt SAVM888 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2488 L=500e-9 W=3e-6
m2 net19 bl 0 0 N888 L=500e-9 W=3e-6
.ends SAVM888

.subckt SAVM889 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2489 L=500e-9 W=3e-6
m2 net19 bl 0 0 N889 L=500e-9 W=3e-6
.ends SAVM889

.subckt SAVM890 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2490 L=500e-9 W=3e-6
m2 net19 bl 0 0 N890 L=500e-9 W=3e-6
.ends SAVM890

.subckt SAVM891 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2491 L=500e-9 W=3e-6
m2 net19 bl 0 0 N891 L=500e-9 W=3e-6
.ends SAVM891

.subckt SAVM892 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2492 L=500e-9 W=3e-6
m2 net19 bl 0 0 N892 L=500e-9 W=3e-6
.ends SAVM892

.subckt SAVM893 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2493 L=500e-9 W=3e-6
m2 net19 bl 0 0 N893 L=500e-9 W=3e-6
.ends SAVM893

.subckt SAVM894 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2494 L=500e-9 W=3e-6
m2 net19 bl 0 0 N894 L=500e-9 W=3e-6
.ends SAVM894

.subckt SAVM895 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2495 L=500e-9 W=3e-6
m2 net19 bl 0 0 N895 L=500e-9 W=3e-6
.ends SAVM895

.subckt SAVM896 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2496 L=500e-9 W=3e-6
m2 net19 bl 0 0 N896 L=500e-9 W=3e-6
.ends SAVM896

.subckt SAVM897 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2497 L=500e-9 W=3e-6
m2 net19 bl 0 0 N897 L=500e-9 W=3e-6
.ends SAVM897

.subckt SAVM898 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2498 L=500e-9 W=3e-6
m2 net19 bl 0 0 N898 L=500e-9 W=3e-6
.ends SAVM898

.subckt SAVM899 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2499 L=500e-9 W=3e-6
m2 net19 bl 0 0 N899 L=500e-9 W=3e-6
.ends SAVM899

.subckt SAVM900 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2500 L=500e-9 W=3e-6
m2 net19 bl 0 0 N900 L=500e-9 W=3e-6
.ends SAVM900

.subckt SAVM901 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2501 L=500e-9 W=3e-6
m2 net19 bl 0 0 N901 L=500e-9 W=3e-6
.ends SAVM901

.subckt SAVM902 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2502 L=500e-9 W=3e-6
m2 net19 bl 0 0 N902 L=500e-9 W=3e-6
.ends SAVM902

.subckt SAVM903 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2503 L=500e-9 W=3e-6
m2 net19 bl 0 0 N903 L=500e-9 W=3e-6
.ends SAVM903

.subckt SAVM904 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2504 L=500e-9 W=3e-6
m2 net19 bl 0 0 N904 L=500e-9 W=3e-6
.ends SAVM904

.subckt SAVM905 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2505 L=500e-9 W=3e-6
m2 net19 bl 0 0 N905 L=500e-9 W=3e-6
.ends SAVM905

.subckt SAVM906 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2506 L=500e-9 W=3e-6
m2 net19 bl 0 0 N906 L=500e-9 W=3e-6
.ends SAVM906

.subckt SAVM907 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2507 L=500e-9 W=3e-6
m2 net19 bl 0 0 N907 L=500e-9 W=3e-6
.ends SAVM907

.subckt SAVM908 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2508 L=500e-9 W=3e-6
m2 net19 bl 0 0 N908 L=500e-9 W=3e-6
.ends SAVM908

.subckt SAVM909 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2509 L=500e-9 W=3e-6
m2 net19 bl 0 0 N909 L=500e-9 W=3e-6
.ends SAVM909

.subckt SAVM910 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2510 L=500e-9 W=3e-6
m2 net19 bl 0 0 N910 L=500e-9 W=3e-6
.ends SAVM910

.subckt SAVM911 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2511 L=500e-9 W=3e-6
m2 net19 bl 0 0 N911 L=500e-9 W=3e-6
.ends SAVM911

.subckt SAVM912 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2512 L=500e-9 W=3e-6
m2 net19 bl 0 0 N912 L=500e-9 W=3e-6
.ends SAVM912

.subckt SAVM913 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2513 L=500e-9 W=3e-6
m2 net19 bl 0 0 N913 L=500e-9 W=3e-6
.ends SAVM913

.subckt SAVM914 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2514 L=500e-9 W=3e-6
m2 net19 bl 0 0 N914 L=500e-9 W=3e-6
.ends SAVM914

.subckt SAVM915 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2515 L=500e-9 W=3e-6
m2 net19 bl 0 0 N915 L=500e-9 W=3e-6
.ends SAVM915

.subckt SAVM916 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2516 L=500e-9 W=3e-6
m2 net19 bl 0 0 N916 L=500e-9 W=3e-6
.ends SAVM916

.subckt SAVM917 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2517 L=500e-9 W=3e-6
m2 net19 bl 0 0 N917 L=500e-9 W=3e-6
.ends SAVM917

.subckt SAVM918 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2518 L=500e-9 W=3e-6
m2 net19 bl 0 0 N918 L=500e-9 W=3e-6
.ends SAVM918

.subckt SAVM919 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2519 L=500e-9 W=3e-6
m2 net19 bl 0 0 N919 L=500e-9 W=3e-6
.ends SAVM919

.subckt SAVM920 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2520 L=500e-9 W=3e-6
m2 net19 bl 0 0 N920 L=500e-9 W=3e-6
.ends SAVM920

.subckt SAVM921 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2521 L=500e-9 W=3e-6
m2 net19 bl 0 0 N921 L=500e-9 W=3e-6
.ends SAVM921

.subckt SAVM922 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2522 L=500e-9 W=3e-6
m2 net19 bl 0 0 N922 L=500e-9 W=3e-6
.ends SAVM922

.subckt SAVM923 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2523 L=500e-9 W=3e-6
m2 net19 bl 0 0 N923 L=500e-9 W=3e-6
.ends SAVM923

.subckt SAVM924 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2524 L=500e-9 W=3e-6
m2 net19 bl 0 0 N924 L=500e-9 W=3e-6
.ends SAVM924

.subckt SAVM925 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2525 L=500e-9 W=3e-6
m2 net19 bl 0 0 N925 L=500e-9 W=3e-6
.ends SAVM925

.subckt SAVM926 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2526 L=500e-9 W=3e-6
m2 net19 bl 0 0 N926 L=500e-9 W=3e-6
.ends SAVM926

.subckt SAVM927 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2527 L=500e-9 W=3e-6
m2 net19 bl 0 0 N927 L=500e-9 W=3e-6
.ends SAVM927

.subckt SAVM928 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2528 L=500e-9 W=3e-6
m2 net19 bl 0 0 N928 L=500e-9 W=3e-6
.ends SAVM928

.subckt SAVM929 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2529 L=500e-9 W=3e-6
m2 net19 bl 0 0 N929 L=500e-9 W=3e-6
.ends SAVM929

.subckt SAVM930 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2530 L=500e-9 W=3e-6
m2 net19 bl 0 0 N930 L=500e-9 W=3e-6
.ends SAVM930

.subckt SAVM931 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2531 L=500e-9 W=3e-6
m2 net19 bl 0 0 N931 L=500e-9 W=3e-6
.ends SAVM931

.subckt SAVM932 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2532 L=500e-9 W=3e-6
m2 net19 bl 0 0 N932 L=500e-9 W=3e-6
.ends SAVM932

.subckt SAVM933 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2533 L=500e-9 W=3e-6
m2 net19 bl 0 0 N933 L=500e-9 W=3e-6
.ends SAVM933

.subckt SAVM934 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2534 L=500e-9 W=3e-6
m2 net19 bl 0 0 N934 L=500e-9 W=3e-6
.ends SAVM934

.subckt SAVM935 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2535 L=500e-9 W=3e-6
m2 net19 bl 0 0 N935 L=500e-9 W=3e-6
.ends SAVM935

.subckt SAVM936 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2536 L=500e-9 W=3e-6
m2 net19 bl 0 0 N936 L=500e-9 W=3e-6
.ends SAVM936

.subckt SAVM937 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2537 L=500e-9 W=3e-6
m2 net19 bl 0 0 N937 L=500e-9 W=3e-6
.ends SAVM937

.subckt SAVM938 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2538 L=500e-9 W=3e-6
m2 net19 bl 0 0 N938 L=500e-9 W=3e-6
.ends SAVM938

.subckt SAVM939 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2539 L=500e-9 W=3e-6
m2 net19 bl 0 0 N939 L=500e-9 W=3e-6
.ends SAVM939

.subckt SAVM940 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2540 L=500e-9 W=3e-6
m2 net19 bl 0 0 N940 L=500e-9 W=3e-6
.ends SAVM940

.subckt SAVM941 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2541 L=500e-9 W=3e-6
m2 net19 bl 0 0 N941 L=500e-9 W=3e-6
.ends SAVM941

.subckt SAVM942 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2542 L=500e-9 W=3e-6
m2 net19 bl 0 0 N942 L=500e-9 W=3e-6
.ends SAVM942

.subckt SAVM943 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2543 L=500e-9 W=3e-6
m2 net19 bl 0 0 N943 L=500e-9 W=3e-6
.ends SAVM943

.subckt SAVM944 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2544 L=500e-9 W=3e-6
m2 net19 bl 0 0 N944 L=500e-9 W=3e-6
.ends SAVM944

.subckt SAVM945 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2545 L=500e-9 W=3e-6
m2 net19 bl 0 0 N945 L=500e-9 W=3e-6
.ends SAVM945

.subckt SAVM946 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2546 L=500e-9 W=3e-6
m2 net19 bl 0 0 N946 L=500e-9 W=3e-6
.ends SAVM946

.subckt SAVM947 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2547 L=500e-9 W=3e-6
m2 net19 bl 0 0 N947 L=500e-9 W=3e-6
.ends SAVM947

.subckt SAVM948 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2548 L=500e-9 W=3e-6
m2 net19 bl 0 0 N948 L=500e-9 W=3e-6
.ends SAVM948

.subckt SAVM949 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2549 L=500e-9 W=3e-6
m2 net19 bl 0 0 N949 L=500e-9 W=3e-6
.ends SAVM949

.subckt SAVM950 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2550 L=500e-9 W=3e-6
m2 net19 bl 0 0 N950 L=500e-9 W=3e-6
.ends SAVM950

.subckt SAVM951 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2551 L=500e-9 W=3e-6
m2 net19 bl 0 0 N951 L=500e-9 W=3e-6
.ends SAVM951

.subckt SAVM952 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2552 L=500e-9 W=3e-6
m2 net19 bl 0 0 N952 L=500e-9 W=3e-6
.ends SAVM952

.subckt SAVM953 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2553 L=500e-9 W=3e-6
m2 net19 bl 0 0 N953 L=500e-9 W=3e-6
.ends SAVM953

.subckt SAVM954 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2554 L=500e-9 W=3e-6
m2 net19 bl 0 0 N954 L=500e-9 W=3e-6
.ends SAVM954

.subckt SAVM955 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2555 L=500e-9 W=3e-6
m2 net19 bl 0 0 N955 L=500e-9 W=3e-6
.ends SAVM955

.subckt SAVM956 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2556 L=500e-9 W=3e-6
m2 net19 bl 0 0 N956 L=500e-9 W=3e-6
.ends SAVM956

.subckt SAVM957 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2557 L=500e-9 W=3e-6
m2 net19 bl 0 0 N957 L=500e-9 W=3e-6
.ends SAVM957

.subckt SAVM958 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2558 L=500e-9 W=3e-6
m2 net19 bl 0 0 N958 L=500e-9 W=3e-6
.ends SAVM958

.subckt SAVM959 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2559 L=500e-9 W=3e-6
m2 net19 bl 0 0 N959 L=500e-9 W=3e-6
.ends SAVM959

.subckt SAVM960 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2560 L=500e-9 W=3e-6
m2 net19 bl 0 0 N960 L=500e-9 W=3e-6
.ends SAVM960

.subckt SAVM961 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2561 L=500e-9 W=3e-6
m2 net19 bl 0 0 N961 L=500e-9 W=3e-6
.ends SAVM961

.subckt SAVM962 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2562 L=500e-9 W=3e-6
m2 net19 bl 0 0 N962 L=500e-9 W=3e-6
.ends SAVM962

.subckt SAVM963 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2563 L=500e-9 W=3e-6
m2 net19 bl 0 0 N963 L=500e-9 W=3e-6
.ends SAVM963

.subckt SAVM964 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2564 L=500e-9 W=3e-6
m2 net19 bl 0 0 N964 L=500e-9 W=3e-6
.ends SAVM964

.subckt SAVM965 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2565 L=500e-9 W=3e-6
m2 net19 bl 0 0 N965 L=500e-9 W=3e-6
.ends SAVM965

.subckt SAVM966 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2566 L=500e-9 W=3e-6
m2 net19 bl 0 0 N966 L=500e-9 W=3e-6
.ends SAVM966

.subckt SAVM967 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2567 L=500e-9 W=3e-6
m2 net19 bl 0 0 N967 L=500e-9 W=3e-6
.ends SAVM967

.subckt SAVM968 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2568 L=500e-9 W=3e-6
m2 net19 bl 0 0 N968 L=500e-9 W=3e-6
.ends SAVM968

.subckt SAVM969 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2569 L=500e-9 W=3e-6
m2 net19 bl 0 0 N969 L=500e-9 W=3e-6
.ends SAVM969

.subckt SAVM970 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2570 L=500e-9 W=3e-6
m2 net19 bl 0 0 N970 L=500e-9 W=3e-6
.ends SAVM970

.subckt SAVM971 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2571 L=500e-9 W=3e-6
m2 net19 bl 0 0 N971 L=500e-9 W=3e-6
.ends SAVM971

.subckt SAVM972 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2572 L=500e-9 W=3e-6
m2 net19 bl 0 0 N972 L=500e-9 W=3e-6
.ends SAVM972

.subckt SAVM973 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2573 L=500e-9 W=3e-6
m2 net19 bl 0 0 N973 L=500e-9 W=3e-6
.ends SAVM973

.subckt SAVM974 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2574 L=500e-9 W=3e-6
m2 net19 bl 0 0 N974 L=500e-9 W=3e-6
.ends SAVM974

.subckt SAVM975 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2575 L=500e-9 W=3e-6
m2 net19 bl 0 0 N975 L=500e-9 W=3e-6
.ends SAVM975

.subckt SAVM976 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2576 L=500e-9 W=3e-6
m2 net19 bl 0 0 N976 L=500e-9 W=3e-6
.ends SAVM976

.subckt SAVM977 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2577 L=500e-9 W=3e-6
m2 net19 bl 0 0 N977 L=500e-9 W=3e-6
.ends SAVM977

.subckt SAVM978 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2578 L=500e-9 W=3e-6
m2 net19 bl 0 0 N978 L=500e-9 W=3e-6
.ends SAVM978

.subckt SAVM979 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2579 L=500e-9 W=3e-6
m2 net19 bl 0 0 N979 L=500e-9 W=3e-6
.ends SAVM979

.subckt SAVM980 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2580 L=500e-9 W=3e-6
m2 net19 bl 0 0 N980 L=500e-9 W=3e-6
.ends SAVM980

.subckt SAVM981 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2581 L=500e-9 W=3e-6
m2 net19 bl 0 0 N981 L=500e-9 W=3e-6
.ends SAVM981

.subckt SAVM982 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2582 L=500e-9 W=3e-6
m2 net19 bl 0 0 N982 L=500e-9 W=3e-6
.ends SAVM982

.subckt SAVM983 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2583 L=500e-9 W=3e-6
m2 net19 bl 0 0 N983 L=500e-9 W=3e-6
.ends SAVM983

.subckt SAVM984 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2584 L=500e-9 W=3e-6
m2 net19 bl 0 0 N984 L=500e-9 W=3e-6
.ends SAVM984

.subckt SAVM985 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2585 L=500e-9 W=3e-6
m2 net19 bl 0 0 N985 L=500e-9 W=3e-6
.ends SAVM985

.subckt SAVM986 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2586 L=500e-9 W=3e-6
m2 net19 bl 0 0 N986 L=500e-9 W=3e-6
.ends SAVM986

.subckt SAVM987 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2587 L=500e-9 W=3e-6
m2 net19 bl 0 0 N987 L=500e-9 W=3e-6
.ends SAVM987

.subckt SAVM988 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2588 L=500e-9 W=3e-6
m2 net19 bl 0 0 N988 L=500e-9 W=3e-6
.ends SAVM988

.subckt SAVM989 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2589 L=500e-9 W=3e-6
m2 net19 bl 0 0 N989 L=500e-9 W=3e-6
.ends SAVM989

.subckt SAVM990 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2590 L=500e-9 W=3e-6
m2 net19 bl 0 0 N990 L=500e-9 W=3e-6
.ends SAVM990

.subckt SAVM991 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2591 L=500e-9 W=3e-6
m2 net19 bl 0 0 N991 L=500e-9 W=3e-6
.ends SAVM991

.subckt SAVM992 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2592 L=500e-9 W=3e-6
m2 net19 bl 0 0 N992 L=500e-9 W=3e-6
.ends SAVM992

.subckt SAVM993 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2593 L=500e-9 W=3e-6
m2 net19 bl 0 0 N993 L=500e-9 W=3e-6
.ends SAVM993

.subckt SAVM994 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2594 L=500e-9 W=3e-6
m2 net19 bl 0 0 N994 L=500e-9 W=3e-6
.ends SAVM994

.subckt SAVM995 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2595 L=500e-9 W=3e-6
m2 net19 bl 0 0 N995 L=500e-9 W=3e-6
.ends SAVM995

.subckt SAVM996 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2596 L=500e-9 W=3e-6
m2 net19 bl 0 0 N996 L=500e-9 W=3e-6
.ends SAVM996

.subckt SAVM997 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2597 L=500e-9 W=3e-6
m2 net19 bl 0 0 N997 L=500e-9 W=3e-6
.ends SAVM997

.subckt SAVM998 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2598 L=500e-9 W=3e-6
m2 net19 bl 0 0 N998 L=500e-9 W=3e-6
.ends SAVM998

.subckt SAVM999 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2599 L=500e-9 W=3e-6
m2 net19 bl 0 0 N999 L=500e-9 W=3e-6
.ends SAVM999

.subckt SAVM1000 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2600 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1000 L=500e-9 W=3e-6
.ends SAVM1000

.subckt SAVM1001 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2601 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1001 L=500e-9 W=3e-6
.ends SAVM1001

.subckt SAVM1002 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2602 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1002 L=500e-9 W=3e-6
.ends SAVM1002

.subckt SAVM1003 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2603 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1003 L=500e-9 W=3e-6
.ends SAVM1003

.subckt SAVM1004 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2604 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1004 L=500e-9 W=3e-6
.ends SAVM1004

.subckt SAVM1005 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2605 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1005 L=500e-9 W=3e-6
.ends SAVM1005

.subckt SAVM1006 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2606 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1006 L=500e-9 W=3e-6
.ends SAVM1006

.subckt SAVM1007 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2607 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1007 L=500e-9 W=3e-6
.ends SAVM1007

.subckt SAVM1008 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2608 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1008 L=500e-9 W=3e-6
.ends SAVM1008

.subckt SAVM1009 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2609 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1009 L=500e-9 W=3e-6
.ends SAVM1009

.subckt SAVM1010 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2610 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1010 L=500e-9 W=3e-6
.ends SAVM1010

.subckt SAVM1011 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2611 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1011 L=500e-9 W=3e-6
.ends SAVM1011

.subckt SAVM1012 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2612 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1012 L=500e-9 W=3e-6
.ends SAVM1012

.subckt SAVM1013 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2613 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1013 L=500e-9 W=3e-6
.ends SAVM1013

.subckt SAVM1014 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2614 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1014 L=500e-9 W=3e-6
.ends SAVM1014

.subckt SAVM1015 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2615 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1015 L=500e-9 W=3e-6
.ends SAVM1015

.subckt SAVM1016 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2616 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1016 L=500e-9 W=3e-6
.ends SAVM1016

.subckt SAVM1017 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2617 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1017 L=500e-9 W=3e-6
.ends SAVM1017

.subckt SAVM1018 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2618 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1018 L=500e-9 W=3e-6
.ends SAVM1018

.subckt SAVM1019 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2619 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1019 L=500e-9 W=3e-6
.ends SAVM1019

.subckt SAVM1020 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2620 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1020 L=500e-9 W=3e-6
.ends SAVM1020

.subckt SAVM1021 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2621 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1021 L=500e-9 W=3e-6
.ends SAVM1021

.subckt SAVM1022 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2622 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1022 L=500e-9 W=3e-6
.ends SAVM1022

.subckt SAVM1023 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2623 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1023 L=500e-9 W=3e-6
.ends SAVM1023

.subckt SAVM1024 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2624 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1024 L=500e-9 W=3e-6
.ends SAVM1024

.subckt SAVM1025 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2625 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1025 L=500e-9 W=3e-6
.ends SAVM1025

.subckt SAVM1026 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2626 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1026 L=500e-9 W=3e-6
.ends SAVM1026

.subckt SAVM1027 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2627 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1027 L=500e-9 W=3e-6
.ends SAVM1027

.subckt SAVM1028 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2628 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1028 L=500e-9 W=3e-6
.ends SAVM1028

.subckt SAVM1029 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2629 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1029 L=500e-9 W=3e-6
.ends SAVM1029

.subckt SAVM1030 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2630 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1030 L=500e-9 W=3e-6
.ends SAVM1030

.subckt SAVM1031 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2631 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1031 L=500e-9 W=3e-6
.ends SAVM1031

.subckt SAVM1032 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2632 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1032 L=500e-9 W=3e-6
.ends SAVM1032

.subckt SAVM1033 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2633 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1033 L=500e-9 W=3e-6
.ends SAVM1033

.subckt SAVM1034 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2634 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1034 L=500e-9 W=3e-6
.ends SAVM1034

.subckt SAVM1035 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2635 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1035 L=500e-9 W=3e-6
.ends SAVM1035

.subckt SAVM1036 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2636 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1036 L=500e-9 W=3e-6
.ends SAVM1036

.subckt SAVM1037 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2637 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1037 L=500e-9 W=3e-6
.ends SAVM1037

.subckt SAVM1038 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2638 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1038 L=500e-9 W=3e-6
.ends SAVM1038

.subckt SAVM1039 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2639 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1039 L=500e-9 W=3e-6
.ends SAVM1039

.subckt SAVM1040 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2640 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1040 L=500e-9 W=3e-6
.ends SAVM1040

.subckt SAVM1041 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2641 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1041 L=500e-9 W=3e-6
.ends SAVM1041

.subckt SAVM1042 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2642 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1042 L=500e-9 W=3e-6
.ends SAVM1042

.subckt SAVM1043 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2643 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1043 L=500e-9 W=3e-6
.ends SAVM1043

.subckt SAVM1044 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2644 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1044 L=500e-9 W=3e-6
.ends SAVM1044

.subckt SAVM1045 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2645 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1045 L=500e-9 W=3e-6
.ends SAVM1045

.subckt SAVM1046 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2646 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1046 L=500e-9 W=3e-6
.ends SAVM1046

.subckt SAVM1047 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2647 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1047 L=500e-9 W=3e-6
.ends SAVM1047

.subckt SAVM1048 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2648 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1048 L=500e-9 W=3e-6
.ends SAVM1048

.subckt SAVM1049 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2649 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1049 L=500e-9 W=3e-6
.ends SAVM1049

.subckt SAVM1050 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2650 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1050 L=500e-9 W=3e-6
.ends SAVM1050

.subckt SAVM1051 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2651 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1051 L=500e-9 W=3e-6
.ends SAVM1051

.subckt SAVM1052 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2652 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1052 L=500e-9 W=3e-6
.ends SAVM1052

.subckt SAVM1053 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2653 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1053 L=500e-9 W=3e-6
.ends SAVM1053

.subckt SAVM1054 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2654 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1054 L=500e-9 W=3e-6
.ends SAVM1054

.subckt SAVM1055 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2655 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1055 L=500e-9 W=3e-6
.ends SAVM1055

.subckt SAVM1056 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2656 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1056 L=500e-9 W=3e-6
.ends SAVM1056

.subckt SAVM1057 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2657 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1057 L=500e-9 W=3e-6
.ends SAVM1057

.subckt SAVM1058 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2658 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1058 L=500e-9 W=3e-6
.ends SAVM1058

.subckt SAVM1059 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2659 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1059 L=500e-9 W=3e-6
.ends SAVM1059

.subckt SAVM1060 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2660 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1060 L=500e-9 W=3e-6
.ends SAVM1060

.subckt SAVM1061 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2661 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1061 L=500e-9 W=3e-6
.ends SAVM1061

.subckt SAVM1062 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2662 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1062 L=500e-9 W=3e-6
.ends SAVM1062

.subckt SAVM1063 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2663 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1063 L=500e-9 W=3e-6
.ends SAVM1063

.subckt SAVM1064 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2664 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1064 L=500e-9 W=3e-6
.ends SAVM1064

.subckt SAVM1065 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2665 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1065 L=500e-9 W=3e-6
.ends SAVM1065

.subckt SAVM1066 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2666 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1066 L=500e-9 W=3e-6
.ends SAVM1066

.subckt SAVM1067 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2667 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1067 L=500e-9 W=3e-6
.ends SAVM1067

.subckt SAVM1068 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2668 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1068 L=500e-9 W=3e-6
.ends SAVM1068

.subckt SAVM1069 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2669 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1069 L=500e-9 W=3e-6
.ends SAVM1069

.subckt SAVM1070 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2670 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1070 L=500e-9 W=3e-6
.ends SAVM1070

.subckt SAVM1071 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2671 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1071 L=500e-9 W=3e-6
.ends SAVM1071

.subckt SAVM1072 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2672 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1072 L=500e-9 W=3e-6
.ends SAVM1072

.subckt SAVM1073 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2673 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1073 L=500e-9 W=3e-6
.ends SAVM1073

.subckt SAVM1074 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2674 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1074 L=500e-9 W=3e-6
.ends SAVM1074

.subckt SAVM1075 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2675 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1075 L=500e-9 W=3e-6
.ends SAVM1075

.subckt SAVM1076 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2676 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1076 L=500e-9 W=3e-6
.ends SAVM1076

.subckt SAVM1077 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2677 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1077 L=500e-9 W=3e-6
.ends SAVM1077

.subckt SAVM1078 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2678 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1078 L=500e-9 W=3e-6
.ends SAVM1078

.subckt SAVM1079 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2679 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1079 L=500e-9 W=3e-6
.ends SAVM1079

.subckt SAVM1080 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2680 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1080 L=500e-9 W=3e-6
.ends SAVM1080

.subckt SAVM1081 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2681 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1081 L=500e-9 W=3e-6
.ends SAVM1081

.subckt SAVM1082 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2682 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1082 L=500e-9 W=3e-6
.ends SAVM1082

.subckt SAVM1083 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2683 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1083 L=500e-9 W=3e-6
.ends SAVM1083

.subckt SAVM1084 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2684 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1084 L=500e-9 W=3e-6
.ends SAVM1084

.subckt SAVM1085 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2685 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1085 L=500e-9 W=3e-6
.ends SAVM1085

.subckt SAVM1086 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2686 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1086 L=500e-9 W=3e-6
.ends SAVM1086

.subckt SAVM1087 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2687 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1087 L=500e-9 W=3e-6
.ends SAVM1087

.subckt SAVM1088 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2688 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1088 L=500e-9 W=3e-6
.ends SAVM1088

.subckt SAVM1089 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2689 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1089 L=500e-9 W=3e-6
.ends SAVM1089

.subckt SAVM1090 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2690 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1090 L=500e-9 W=3e-6
.ends SAVM1090

.subckt SAVM1091 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2691 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1091 L=500e-9 W=3e-6
.ends SAVM1091

.subckt SAVM1092 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2692 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1092 L=500e-9 W=3e-6
.ends SAVM1092

.subckt SAVM1093 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2693 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1093 L=500e-9 W=3e-6
.ends SAVM1093

.subckt SAVM1094 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2694 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1094 L=500e-9 W=3e-6
.ends SAVM1094

.subckt SAVM1095 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2695 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1095 L=500e-9 W=3e-6
.ends SAVM1095

.subckt SAVM1096 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2696 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1096 L=500e-9 W=3e-6
.ends SAVM1096

.subckt SAVM1097 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2697 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1097 L=500e-9 W=3e-6
.ends SAVM1097

.subckt SAVM1098 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2698 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1098 L=500e-9 W=3e-6
.ends SAVM1098

.subckt SAVM1099 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2699 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1099 L=500e-9 W=3e-6
.ends SAVM1099

.subckt SAVM1100 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2700 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1100 L=500e-9 W=3e-6
.ends SAVM1100

.subckt SAVM1101 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2701 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1101 L=500e-9 W=3e-6
.ends SAVM1101

.subckt SAVM1102 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2702 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1102 L=500e-9 W=3e-6
.ends SAVM1102

.subckt SAVM1103 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2703 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1103 L=500e-9 W=3e-6
.ends SAVM1103

.subckt SAVM1104 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2704 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1104 L=500e-9 W=3e-6
.ends SAVM1104

.subckt SAVM1105 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2705 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1105 L=500e-9 W=3e-6
.ends SAVM1105

.subckt SAVM1106 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2706 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1106 L=500e-9 W=3e-6
.ends SAVM1106

.subckt SAVM1107 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2707 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1107 L=500e-9 W=3e-6
.ends SAVM1107

.subckt SAVM1108 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2708 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1108 L=500e-9 W=3e-6
.ends SAVM1108

.subckt SAVM1109 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2709 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1109 L=500e-9 W=3e-6
.ends SAVM1109

.subckt SAVM1110 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2710 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1110 L=500e-9 W=3e-6
.ends SAVM1110

.subckt SAVM1111 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2711 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1111 L=500e-9 W=3e-6
.ends SAVM1111

.subckt SAVM1112 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2712 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1112 L=500e-9 W=3e-6
.ends SAVM1112

.subckt SAVM1113 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2713 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1113 L=500e-9 W=3e-6
.ends SAVM1113

.subckt SAVM1114 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2714 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1114 L=500e-9 W=3e-6
.ends SAVM1114

.subckt SAVM1115 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2715 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1115 L=500e-9 W=3e-6
.ends SAVM1115

.subckt SAVM1116 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2716 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1116 L=500e-9 W=3e-6
.ends SAVM1116

.subckt SAVM1117 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2717 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1117 L=500e-9 W=3e-6
.ends SAVM1117

.subckt SAVM1118 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2718 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1118 L=500e-9 W=3e-6
.ends SAVM1118

.subckt SAVM1119 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2719 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1119 L=500e-9 W=3e-6
.ends SAVM1119

.subckt SAVM1120 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2720 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1120 L=500e-9 W=3e-6
.ends SAVM1120

.subckt SAVM1121 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2721 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1121 L=500e-9 W=3e-6
.ends SAVM1121

.subckt SAVM1122 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2722 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1122 L=500e-9 W=3e-6
.ends SAVM1122

.subckt SAVM1123 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2723 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1123 L=500e-9 W=3e-6
.ends SAVM1123

.subckt SAVM1124 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2724 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1124 L=500e-9 W=3e-6
.ends SAVM1124

.subckt SAVM1125 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2725 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1125 L=500e-9 W=3e-6
.ends SAVM1125

.subckt SAVM1126 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2726 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1126 L=500e-9 W=3e-6
.ends SAVM1126

.subckt SAVM1127 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2727 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1127 L=500e-9 W=3e-6
.ends SAVM1127

.subckt SAVM1128 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2728 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1128 L=500e-9 W=3e-6
.ends SAVM1128

.subckt SAVM1129 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2729 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1129 L=500e-9 W=3e-6
.ends SAVM1129

.subckt SAVM1130 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2730 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1130 L=500e-9 W=3e-6
.ends SAVM1130

.subckt SAVM1131 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2731 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1131 L=500e-9 W=3e-6
.ends SAVM1131

.subckt SAVM1132 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2732 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1132 L=500e-9 W=3e-6
.ends SAVM1132

.subckt SAVM1133 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2733 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1133 L=500e-9 W=3e-6
.ends SAVM1133

.subckt SAVM1134 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2734 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1134 L=500e-9 W=3e-6
.ends SAVM1134

.subckt SAVM1135 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2735 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1135 L=500e-9 W=3e-6
.ends SAVM1135

.subckt SAVM1136 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2736 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1136 L=500e-9 W=3e-6
.ends SAVM1136

.subckt SAVM1137 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2737 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1137 L=500e-9 W=3e-6
.ends SAVM1137

.subckt SAVM1138 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2738 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1138 L=500e-9 W=3e-6
.ends SAVM1138

.subckt SAVM1139 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2739 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1139 L=500e-9 W=3e-6
.ends SAVM1139

.subckt SAVM1140 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2740 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1140 L=500e-9 W=3e-6
.ends SAVM1140

.subckt SAVM1141 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2741 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1141 L=500e-9 W=3e-6
.ends SAVM1141

.subckt SAVM1142 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2742 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1142 L=500e-9 W=3e-6
.ends SAVM1142

.subckt SAVM1143 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2743 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1143 L=500e-9 W=3e-6
.ends SAVM1143

.subckt SAVM1144 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2744 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1144 L=500e-9 W=3e-6
.ends SAVM1144

.subckt SAVM1145 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2745 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1145 L=500e-9 W=3e-6
.ends SAVM1145

.subckt SAVM1146 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2746 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1146 L=500e-9 W=3e-6
.ends SAVM1146

.subckt SAVM1147 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2747 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1147 L=500e-9 W=3e-6
.ends SAVM1147

.subckt SAVM1148 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2748 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1148 L=500e-9 W=3e-6
.ends SAVM1148

.subckt SAVM1149 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2749 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1149 L=500e-9 W=3e-6
.ends SAVM1149

.subckt SAVM1150 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2750 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1150 L=500e-9 W=3e-6
.ends SAVM1150

.subckt SAVM1151 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2751 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1151 L=500e-9 W=3e-6
.ends SAVM1151

.subckt SAVM1152 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2752 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1152 L=500e-9 W=3e-6
.ends SAVM1152

.subckt SAVM1153 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2753 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1153 L=500e-9 W=3e-6
.ends SAVM1153

.subckt SAVM1154 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2754 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1154 L=500e-9 W=3e-6
.ends SAVM1154

.subckt SAVM1155 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2755 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1155 L=500e-9 W=3e-6
.ends SAVM1155

.subckt SAVM1156 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2756 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1156 L=500e-9 W=3e-6
.ends SAVM1156

.subckt SAVM1157 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2757 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1157 L=500e-9 W=3e-6
.ends SAVM1157

.subckt SAVM1158 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2758 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1158 L=500e-9 W=3e-6
.ends SAVM1158

.subckt SAVM1159 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2759 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1159 L=500e-9 W=3e-6
.ends SAVM1159

.subckt SAVM1160 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2760 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1160 L=500e-9 W=3e-6
.ends SAVM1160

.subckt SAVM1161 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2761 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1161 L=500e-9 W=3e-6
.ends SAVM1161

.subckt SAVM1162 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2762 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1162 L=500e-9 W=3e-6
.ends SAVM1162

.subckt SAVM1163 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2763 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1163 L=500e-9 W=3e-6
.ends SAVM1163

.subckt SAVM1164 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2764 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1164 L=500e-9 W=3e-6
.ends SAVM1164

.subckt SAVM1165 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2765 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1165 L=500e-9 W=3e-6
.ends SAVM1165

.subckt SAVM1166 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2766 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1166 L=500e-9 W=3e-6
.ends SAVM1166

.subckt SAVM1167 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2767 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1167 L=500e-9 W=3e-6
.ends SAVM1167

.subckt SAVM1168 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2768 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1168 L=500e-9 W=3e-6
.ends SAVM1168

.subckt SAVM1169 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2769 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1169 L=500e-9 W=3e-6
.ends SAVM1169

.subckt SAVM1170 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2770 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1170 L=500e-9 W=3e-6
.ends SAVM1170

.subckt SAVM1171 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2771 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1171 L=500e-9 W=3e-6
.ends SAVM1171

.subckt SAVM1172 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2772 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1172 L=500e-9 W=3e-6
.ends SAVM1172

.subckt SAVM1173 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2773 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1173 L=500e-9 W=3e-6
.ends SAVM1173

.subckt SAVM1174 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2774 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1174 L=500e-9 W=3e-6
.ends SAVM1174

.subckt SAVM1175 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2775 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1175 L=500e-9 W=3e-6
.ends SAVM1175

.subckt SAVM1176 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2776 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1176 L=500e-9 W=3e-6
.ends SAVM1176

.subckt SAVM1177 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2777 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1177 L=500e-9 W=3e-6
.ends SAVM1177

.subckt SAVM1178 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2778 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1178 L=500e-9 W=3e-6
.ends SAVM1178

.subckt SAVM1179 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2779 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1179 L=500e-9 W=3e-6
.ends SAVM1179

.subckt SAVM1180 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2780 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1180 L=500e-9 W=3e-6
.ends SAVM1180

.subckt SAVM1181 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2781 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1181 L=500e-9 W=3e-6
.ends SAVM1181

.subckt SAVM1182 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2782 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1182 L=500e-9 W=3e-6
.ends SAVM1182

.subckt SAVM1183 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2783 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1183 L=500e-9 W=3e-6
.ends SAVM1183

.subckt SAVM1184 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2784 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1184 L=500e-9 W=3e-6
.ends SAVM1184

.subckt SAVM1185 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2785 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1185 L=500e-9 W=3e-6
.ends SAVM1185

.subckt SAVM1186 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2786 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1186 L=500e-9 W=3e-6
.ends SAVM1186

.subckt SAVM1187 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2787 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1187 L=500e-9 W=3e-6
.ends SAVM1187

.subckt SAVM1188 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2788 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1188 L=500e-9 W=3e-6
.ends SAVM1188

.subckt SAVM1189 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2789 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1189 L=500e-9 W=3e-6
.ends SAVM1189

.subckt SAVM1190 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2790 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1190 L=500e-9 W=3e-6
.ends SAVM1190

.subckt SAVM1191 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2791 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1191 L=500e-9 W=3e-6
.ends SAVM1191

.subckt SAVM1192 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2792 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1192 L=500e-9 W=3e-6
.ends SAVM1192

.subckt SAVM1193 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2793 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1193 L=500e-9 W=3e-6
.ends SAVM1193

.subckt SAVM1194 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2794 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1194 L=500e-9 W=3e-6
.ends SAVM1194

.subckt SAVM1195 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2795 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1195 L=500e-9 W=3e-6
.ends SAVM1195

.subckt SAVM1196 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2796 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1196 L=500e-9 W=3e-6
.ends SAVM1196

.subckt SAVM1197 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2797 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1197 L=500e-9 W=3e-6
.ends SAVM1197

.subckt SAVM1198 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2798 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1198 L=500e-9 W=3e-6
.ends SAVM1198

.subckt SAVM1199 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2799 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1199 L=500e-9 W=3e-6
.ends SAVM1199

.subckt SAVM1200 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2800 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1200 L=500e-9 W=3e-6
.ends SAVM1200

.subckt SAVM1201 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2801 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1201 L=500e-9 W=3e-6
.ends SAVM1201

.subckt SAVM1202 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2802 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1202 L=500e-9 W=3e-6
.ends SAVM1202

.subckt SAVM1203 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2803 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1203 L=500e-9 W=3e-6
.ends SAVM1203

.subckt SAVM1204 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2804 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1204 L=500e-9 W=3e-6
.ends SAVM1204

.subckt SAVM1205 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2805 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1205 L=500e-9 W=3e-6
.ends SAVM1205

.subckt SAVM1206 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2806 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1206 L=500e-9 W=3e-6
.ends SAVM1206

.subckt SAVM1207 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2807 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1207 L=500e-9 W=3e-6
.ends SAVM1207

.subckt SAVM1208 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2808 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1208 L=500e-9 W=3e-6
.ends SAVM1208

.subckt SAVM1209 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2809 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1209 L=500e-9 W=3e-6
.ends SAVM1209

.subckt SAVM1210 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2810 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1210 L=500e-9 W=3e-6
.ends SAVM1210

.subckt SAVM1211 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2811 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1211 L=500e-9 W=3e-6
.ends SAVM1211

.subckt SAVM1212 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2812 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1212 L=500e-9 W=3e-6
.ends SAVM1212

.subckt SAVM1213 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2813 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1213 L=500e-9 W=3e-6
.ends SAVM1213

.subckt SAVM1214 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2814 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1214 L=500e-9 W=3e-6
.ends SAVM1214

.subckt SAVM1215 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2815 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1215 L=500e-9 W=3e-6
.ends SAVM1215

.subckt SAVM1216 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2816 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1216 L=500e-9 W=3e-6
.ends SAVM1216

.subckt SAVM1217 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2817 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1217 L=500e-9 W=3e-6
.ends SAVM1217

.subckt SAVM1218 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2818 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1218 L=500e-9 W=3e-6
.ends SAVM1218

.subckt SAVM1219 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2819 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1219 L=500e-9 W=3e-6
.ends SAVM1219

.subckt SAVM1220 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2820 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1220 L=500e-9 W=3e-6
.ends SAVM1220

.subckt SAVM1221 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2821 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1221 L=500e-9 W=3e-6
.ends SAVM1221

.subckt SAVM1222 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2822 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1222 L=500e-9 W=3e-6
.ends SAVM1222

.subckt SAVM1223 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2823 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1223 L=500e-9 W=3e-6
.ends SAVM1223

.subckt SAVM1224 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2824 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1224 L=500e-9 W=3e-6
.ends SAVM1224

.subckt SAVM1225 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2825 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1225 L=500e-9 W=3e-6
.ends SAVM1225

.subckt SAVM1226 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2826 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1226 L=500e-9 W=3e-6
.ends SAVM1226

.subckt SAVM1227 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2827 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1227 L=500e-9 W=3e-6
.ends SAVM1227

.subckt SAVM1228 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2828 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1228 L=500e-9 W=3e-6
.ends SAVM1228

.subckt SAVM1229 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2829 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1229 L=500e-9 W=3e-6
.ends SAVM1229

.subckt SAVM1230 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2830 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1230 L=500e-9 W=3e-6
.ends SAVM1230

.subckt SAVM1231 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2831 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1231 L=500e-9 W=3e-6
.ends SAVM1231

.subckt SAVM1232 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2832 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1232 L=500e-9 W=3e-6
.ends SAVM1232

.subckt SAVM1233 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2833 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1233 L=500e-9 W=3e-6
.ends SAVM1233

.subckt SAVM1234 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2834 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1234 L=500e-9 W=3e-6
.ends SAVM1234

.subckt SAVM1235 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2835 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1235 L=500e-9 W=3e-6
.ends SAVM1235

.subckt SAVM1236 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2836 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1236 L=500e-9 W=3e-6
.ends SAVM1236

.subckt SAVM1237 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2837 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1237 L=500e-9 W=3e-6
.ends SAVM1237

.subckt SAVM1238 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2838 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1238 L=500e-9 W=3e-6
.ends SAVM1238

.subckt SAVM1239 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2839 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1239 L=500e-9 W=3e-6
.ends SAVM1239

.subckt SAVM1240 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2840 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1240 L=500e-9 W=3e-6
.ends SAVM1240

.subckt SAVM1241 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2841 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1241 L=500e-9 W=3e-6
.ends SAVM1241

.subckt SAVM1242 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2842 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1242 L=500e-9 W=3e-6
.ends SAVM1242

.subckt SAVM1243 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2843 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1243 L=500e-9 W=3e-6
.ends SAVM1243

.subckt SAVM1244 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2844 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1244 L=500e-9 W=3e-6
.ends SAVM1244

.subckt SAVM1245 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2845 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1245 L=500e-9 W=3e-6
.ends SAVM1245

.subckt SAVM1246 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2846 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1246 L=500e-9 W=3e-6
.ends SAVM1246

.subckt SAVM1247 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2847 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1247 L=500e-9 W=3e-6
.ends SAVM1247

.subckt SAVM1248 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2848 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1248 L=500e-9 W=3e-6
.ends SAVM1248

.subckt SAVM1249 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2849 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1249 L=500e-9 W=3e-6
.ends SAVM1249

.subckt SAVM1250 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2850 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1250 L=500e-9 W=3e-6
.ends SAVM1250

.subckt SAVM1251 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2851 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1251 L=500e-9 W=3e-6
.ends SAVM1251

.subckt SAVM1252 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2852 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1252 L=500e-9 W=3e-6
.ends SAVM1252

.subckt SAVM1253 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2853 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1253 L=500e-9 W=3e-6
.ends SAVM1253

.subckt SAVM1254 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2854 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1254 L=500e-9 W=3e-6
.ends SAVM1254

.subckt SAVM1255 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2855 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1255 L=500e-9 W=3e-6
.ends SAVM1255

.subckt SAVM1256 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2856 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1256 L=500e-9 W=3e-6
.ends SAVM1256

.subckt SAVM1257 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2857 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1257 L=500e-9 W=3e-6
.ends SAVM1257

.subckt SAVM1258 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2858 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1258 L=500e-9 W=3e-6
.ends SAVM1258

.subckt SAVM1259 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2859 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1259 L=500e-9 W=3e-6
.ends SAVM1259

.subckt SAVM1260 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2860 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1260 L=500e-9 W=3e-6
.ends SAVM1260

.subckt SAVM1261 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2861 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1261 L=500e-9 W=3e-6
.ends SAVM1261

.subckt SAVM1262 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2862 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1262 L=500e-9 W=3e-6
.ends SAVM1262

.subckt SAVM1263 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2863 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1263 L=500e-9 W=3e-6
.ends SAVM1263

.subckt SAVM1264 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2864 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1264 L=500e-9 W=3e-6
.ends SAVM1264

.subckt SAVM1265 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2865 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1265 L=500e-9 W=3e-6
.ends SAVM1265

.subckt SAVM1266 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2866 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1266 L=500e-9 W=3e-6
.ends SAVM1266

.subckt SAVM1267 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2867 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1267 L=500e-9 W=3e-6
.ends SAVM1267

.subckt SAVM1268 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2868 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1268 L=500e-9 W=3e-6
.ends SAVM1268

.subckt SAVM1269 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2869 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1269 L=500e-9 W=3e-6
.ends SAVM1269

.subckt SAVM1270 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2870 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1270 L=500e-9 W=3e-6
.ends SAVM1270

.subckt SAVM1271 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2871 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1271 L=500e-9 W=3e-6
.ends SAVM1271

.subckt SAVM1272 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2872 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1272 L=500e-9 W=3e-6
.ends SAVM1272

.subckt SAVM1273 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2873 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1273 L=500e-9 W=3e-6
.ends SAVM1273

.subckt SAVM1274 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2874 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1274 L=500e-9 W=3e-6
.ends SAVM1274

.subckt SAVM1275 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2875 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1275 L=500e-9 W=3e-6
.ends SAVM1275

.subckt SAVM1276 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2876 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1276 L=500e-9 W=3e-6
.ends SAVM1276

.subckt SAVM1277 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2877 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1277 L=500e-9 W=3e-6
.ends SAVM1277

.subckt SAVM1278 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2878 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1278 L=500e-9 W=3e-6
.ends SAVM1278

.subckt SAVM1279 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2879 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1279 L=500e-9 W=3e-6
.ends SAVM1279

.subckt SAVM1280 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2880 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1280 L=500e-9 W=3e-6
.ends SAVM1280

.subckt SAVM1281 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2881 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1281 L=500e-9 W=3e-6
.ends SAVM1281

.subckt SAVM1282 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2882 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1282 L=500e-9 W=3e-6
.ends SAVM1282

.subckt SAVM1283 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2883 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1283 L=500e-9 W=3e-6
.ends SAVM1283

.subckt SAVM1284 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2884 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1284 L=500e-9 W=3e-6
.ends SAVM1284

.subckt SAVM1285 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2885 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1285 L=500e-9 W=3e-6
.ends SAVM1285

.subckt SAVM1286 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2886 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1286 L=500e-9 W=3e-6
.ends SAVM1286

.subckt SAVM1287 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2887 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1287 L=500e-9 W=3e-6
.ends SAVM1287

.subckt SAVM1288 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2888 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1288 L=500e-9 W=3e-6
.ends SAVM1288

.subckt SAVM1289 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2889 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1289 L=500e-9 W=3e-6
.ends SAVM1289

.subckt SAVM1290 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2890 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1290 L=500e-9 W=3e-6
.ends SAVM1290

.subckt SAVM1291 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2891 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1291 L=500e-9 W=3e-6
.ends SAVM1291

.subckt SAVM1292 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2892 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1292 L=500e-9 W=3e-6
.ends SAVM1292

.subckt SAVM1293 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2893 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1293 L=500e-9 W=3e-6
.ends SAVM1293

.subckt SAVM1294 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2894 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1294 L=500e-9 W=3e-6
.ends SAVM1294

.subckt SAVM1295 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2895 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1295 L=500e-9 W=3e-6
.ends SAVM1295

.subckt SAVM1296 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2896 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1296 L=500e-9 W=3e-6
.ends SAVM1296

.subckt SAVM1297 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2897 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1297 L=500e-9 W=3e-6
.ends SAVM1297

.subckt SAVM1298 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2898 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1298 L=500e-9 W=3e-6
.ends SAVM1298

.subckt SAVM1299 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2899 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1299 L=500e-9 W=3e-6
.ends SAVM1299

.subckt SAVM1300 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2900 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1300 L=500e-9 W=3e-6
.ends SAVM1300

.subckt SAVM1301 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2901 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1301 L=500e-9 W=3e-6
.ends SAVM1301

.subckt SAVM1302 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2902 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1302 L=500e-9 W=3e-6
.ends SAVM1302

.subckt SAVM1303 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2903 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1303 L=500e-9 W=3e-6
.ends SAVM1303

.subckt SAVM1304 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2904 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1304 L=500e-9 W=3e-6
.ends SAVM1304

.subckt SAVM1305 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2905 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1305 L=500e-9 W=3e-6
.ends SAVM1305

.subckt SAVM1306 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2906 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1306 L=500e-9 W=3e-6
.ends SAVM1306

.subckt SAVM1307 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2907 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1307 L=500e-9 W=3e-6
.ends SAVM1307

.subckt SAVM1308 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2908 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1308 L=500e-9 W=3e-6
.ends SAVM1308

.subckt SAVM1309 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2909 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1309 L=500e-9 W=3e-6
.ends SAVM1309

.subckt SAVM1310 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2910 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1310 L=500e-9 W=3e-6
.ends SAVM1310

.subckt SAVM1311 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2911 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1311 L=500e-9 W=3e-6
.ends SAVM1311

.subckt SAVM1312 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2912 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1312 L=500e-9 W=3e-6
.ends SAVM1312

.subckt SAVM1313 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2913 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1313 L=500e-9 W=3e-6
.ends SAVM1313

.subckt SAVM1314 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2914 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1314 L=500e-9 W=3e-6
.ends SAVM1314

.subckt SAVM1315 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2915 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1315 L=500e-9 W=3e-6
.ends SAVM1315

.subckt SAVM1316 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2916 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1316 L=500e-9 W=3e-6
.ends SAVM1316

.subckt SAVM1317 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2917 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1317 L=500e-9 W=3e-6
.ends SAVM1317

.subckt SAVM1318 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2918 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1318 L=500e-9 W=3e-6
.ends SAVM1318

.subckt SAVM1319 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2919 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1319 L=500e-9 W=3e-6
.ends SAVM1319

.subckt SAVM1320 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2920 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1320 L=500e-9 W=3e-6
.ends SAVM1320

.subckt SAVM1321 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2921 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1321 L=500e-9 W=3e-6
.ends SAVM1321

.subckt SAVM1322 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2922 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1322 L=500e-9 W=3e-6
.ends SAVM1322

.subckt SAVM1323 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2923 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1323 L=500e-9 W=3e-6
.ends SAVM1323

.subckt SAVM1324 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2924 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1324 L=500e-9 W=3e-6
.ends SAVM1324

.subckt SAVM1325 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2925 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1325 L=500e-9 W=3e-6
.ends SAVM1325

.subckt SAVM1326 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2926 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1326 L=500e-9 W=3e-6
.ends SAVM1326

.subckt SAVM1327 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2927 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1327 L=500e-9 W=3e-6
.ends SAVM1327

.subckt SAVM1328 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2928 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1328 L=500e-9 W=3e-6
.ends SAVM1328

.subckt SAVM1329 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2929 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1329 L=500e-9 W=3e-6
.ends SAVM1329

.subckt SAVM1330 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2930 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1330 L=500e-9 W=3e-6
.ends SAVM1330

.subckt SAVM1331 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2931 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1331 L=500e-9 W=3e-6
.ends SAVM1331

.subckt SAVM1332 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2932 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1332 L=500e-9 W=3e-6
.ends SAVM1332

.subckt SAVM1333 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2933 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1333 L=500e-9 W=3e-6
.ends SAVM1333

.subckt SAVM1334 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2934 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1334 L=500e-9 W=3e-6
.ends SAVM1334

.subckt SAVM1335 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2935 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1335 L=500e-9 W=3e-6
.ends SAVM1335

.subckt SAVM1336 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2936 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1336 L=500e-9 W=3e-6
.ends SAVM1336

.subckt SAVM1337 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2937 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1337 L=500e-9 W=3e-6
.ends SAVM1337

.subckt SAVM1338 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2938 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1338 L=500e-9 W=3e-6
.ends SAVM1338

.subckt SAVM1339 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2939 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1339 L=500e-9 W=3e-6
.ends SAVM1339

.subckt SAVM1340 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2940 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1340 L=500e-9 W=3e-6
.ends SAVM1340

.subckt SAVM1341 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2941 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1341 L=500e-9 W=3e-6
.ends SAVM1341

.subckt SAVM1342 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2942 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1342 L=500e-9 W=3e-6
.ends SAVM1342

.subckt SAVM1343 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2943 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1343 L=500e-9 W=3e-6
.ends SAVM1343

.subckt SAVM1344 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2944 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1344 L=500e-9 W=3e-6
.ends SAVM1344

.subckt SAVM1345 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2945 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1345 L=500e-9 W=3e-6
.ends SAVM1345

.subckt SAVM1346 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2946 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1346 L=500e-9 W=3e-6
.ends SAVM1346

.subckt SAVM1347 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2947 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1347 L=500e-9 W=3e-6
.ends SAVM1347

.subckt SAVM1348 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2948 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1348 L=500e-9 W=3e-6
.ends SAVM1348

.subckt SAVM1349 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2949 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1349 L=500e-9 W=3e-6
.ends SAVM1349

.subckt SAVM1350 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2950 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1350 L=500e-9 W=3e-6
.ends SAVM1350

.subckt SAVM1351 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2951 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1351 L=500e-9 W=3e-6
.ends SAVM1351

.subckt SAVM1352 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2952 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1352 L=500e-9 W=3e-6
.ends SAVM1352

.subckt SAVM1353 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2953 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1353 L=500e-9 W=3e-6
.ends SAVM1353

.subckt SAVM1354 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2954 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1354 L=500e-9 W=3e-6
.ends SAVM1354

.subckt SAVM1355 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2955 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1355 L=500e-9 W=3e-6
.ends SAVM1355

.subckt SAVM1356 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2956 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1356 L=500e-9 W=3e-6
.ends SAVM1356

.subckt SAVM1357 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2957 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1357 L=500e-9 W=3e-6
.ends SAVM1357

.subckt SAVM1358 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2958 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1358 L=500e-9 W=3e-6
.ends SAVM1358

.subckt SAVM1359 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2959 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1359 L=500e-9 W=3e-6
.ends SAVM1359

.subckt SAVM1360 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2960 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1360 L=500e-9 W=3e-6
.ends SAVM1360

.subckt SAVM1361 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2961 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1361 L=500e-9 W=3e-6
.ends SAVM1361

.subckt SAVM1362 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2962 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1362 L=500e-9 W=3e-6
.ends SAVM1362

.subckt SAVM1363 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2963 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1363 L=500e-9 W=3e-6
.ends SAVM1363

.subckt SAVM1364 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2964 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1364 L=500e-9 W=3e-6
.ends SAVM1364

.subckt SAVM1365 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2965 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1365 L=500e-9 W=3e-6
.ends SAVM1365

.subckt SAVM1366 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2966 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1366 L=500e-9 W=3e-6
.ends SAVM1366

.subckt SAVM1367 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2967 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1367 L=500e-9 W=3e-6
.ends SAVM1367

.subckt SAVM1368 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2968 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1368 L=500e-9 W=3e-6
.ends SAVM1368

.subckt SAVM1369 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2969 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1369 L=500e-9 W=3e-6
.ends SAVM1369

.subckt SAVM1370 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2970 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1370 L=500e-9 W=3e-6
.ends SAVM1370

.subckt SAVM1371 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2971 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1371 L=500e-9 W=3e-6
.ends SAVM1371

.subckt SAVM1372 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2972 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1372 L=500e-9 W=3e-6
.ends SAVM1372

.subckt SAVM1373 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2973 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1373 L=500e-9 W=3e-6
.ends SAVM1373

.subckt SAVM1374 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2974 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1374 L=500e-9 W=3e-6
.ends SAVM1374

.subckt SAVM1375 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2975 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1375 L=500e-9 W=3e-6
.ends SAVM1375

.subckt SAVM1376 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2976 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1376 L=500e-9 W=3e-6
.ends SAVM1376

.subckt SAVM1377 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2977 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1377 L=500e-9 W=3e-6
.ends SAVM1377

.subckt SAVM1378 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2978 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1378 L=500e-9 W=3e-6
.ends SAVM1378

.subckt SAVM1379 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2979 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1379 L=500e-9 W=3e-6
.ends SAVM1379

.subckt SAVM1380 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2980 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1380 L=500e-9 W=3e-6
.ends SAVM1380

.subckt SAVM1381 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2981 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1381 L=500e-9 W=3e-6
.ends SAVM1381

.subckt SAVM1382 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2982 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1382 L=500e-9 W=3e-6
.ends SAVM1382

.subckt SAVM1383 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2983 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1383 L=500e-9 W=3e-6
.ends SAVM1383

.subckt SAVM1384 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2984 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1384 L=500e-9 W=3e-6
.ends SAVM1384

.subckt SAVM1385 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2985 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1385 L=500e-9 W=3e-6
.ends SAVM1385

.subckt SAVM1386 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2986 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1386 L=500e-9 W=3e-6
.ends SAVM1386

.subckt SAVM1387 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2987 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1387 L=500e-9 W=3e-6
.ends SAVM1387

.subckt SAVM1388 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2988 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1388 L=500e-9 W=3e-6
.ends SAVM1388

.subckt SAVM1389 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2989 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1389 L=500e-9 W=3e-6
.ends SAVM1389

.subckt SAVM1390 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2990 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1390 L=500e-9 W=3e-6
.ends SAVM1390

.subckt SAVM1391 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2991 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1391 L=500e-9 W=3e-6
.ends SAVM1391

.subckt SAVM1392 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2992 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1392 L=500e-9 W=3e-6
.ends SAVM1392

.subckt SAVM1393 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2993 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1393 L=500e-9 W=3e-6
.ends SAVM1393

.subckt SAVM1394 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2994 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1394 L=500e-9 W=3e-6
.ends SAVM1394

.subckt SAVM1395 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2995 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1395 L=500e-9 W=3e-6
.ends SAVM1395

.subckt SAVM1396 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2996 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1396 L=500e-9 W=3e-6
.ends SAVM1396

.subckt SAVM1397 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2997 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1397 L=500e-9 W=3e-6
.ends SAVM1397

.subckt SAVM1398 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2998 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1398 L=500e-9 W=3e-6
.ends SAVM1398

.subckt SAVM1399 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N2999 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1399 L=500e-9 W=3e-6
.ends SAVM1399

.subckt SAVM1400 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3000 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1400 L=500e-9 W=3e-6
.ends SAVM1400

.subckt SAVM1401 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3001 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1401 L=500e-9 W=3e-6
.ends SAVM1401

.subckt SAVM1402 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3002 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1402 L=500e-9 W=3e-6
.ends SAVM1402

.subckt SAVM1403 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3003 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1403 L=500e-9 W=3e-6
.ends SAVM1403

.subckt SAVM1404 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3004 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1404 L=500e-9 W=3e-6
.ends SAVM1404

.subckt SAVM1405 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3005 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1405 L=500e-9 W=3e-6
.ends SAVM1405

.subckt SAVM1406 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3006 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1406 L=500e-9 W=3e-6
.ends SAVM1406

.subckt SAVM1407 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3007 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1407 L=500e-9 W=3e-6
.ends SAVM1407

.subckt SAVM1408 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3008 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1408 L=500e-9 W=3e-6
.ends SAVM1408

.subckt SAVM1409 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3009 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1409 L=500e-9 W=3e-6
.ends SAVM1409

.subckt SAVM1410 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3010 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1410 L=500e-9 W=3e-6
.ends SAVM1410

.subckt SAVM1411 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3011 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1411 L=500e-9 W=3e-6
.ends SAVM1411

.subckt SAVM1412 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3012 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1412 L=500e-9 W=3e-6
.ends SAVM1412

.subckt SAVM1413 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3013 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1413 L=500e-9 W=3e-6
.ends SAVM1413

.subckt SAVM1414 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3014 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1414 L=500e-9 W=3e-6
.ends SAVM1414

.subckt SAVM1415 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3015 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1415 L=500e-9 W=3e-6
.ends SAVM1415

.subckt SAVM1416 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3016 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1416 L=500e-9 W=3e-6
.ends SAVM1416

.subckt SAVM1417 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3017 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1417 L=500e-9 W=3e-6
.ends SAVM1417

.subckt SAVM1418 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3018 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1418 L=500e-9 W=3e-6
.ends SAVM1418

.subckt SAVM1419 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3019 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1419 L=500e-9 W=3e-6
.ends SAVM1419

.subckt SAVM1420 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3020 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1420 L=500e-9 W=3e-6
.ends SAVM1420

.subckt SAVM1421 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3021 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1421 L=500e-9 W=3e-6
.ends SAVM1421

.subckt SAVM1422 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3022 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1422 L=500e-9 W=3e-6
.ends SAVM1422

.subckt SAVM1423 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3023 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1423 L=500e-9 W=3e-6
.ends SAVM1423

.subckt SAVM1424 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3024 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1424 L=500e-9 W=3e-6
.ends SAVM1424

.subckt SAVM1425 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3025 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1425 L=500e-9 W=3e-6
.ends SAVM1425

.subckt SAVM1426 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3026 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1426 L=500e-9 W=3e-6
.ends SAVM1426

.subckt SAVM1427 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3027 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1427 L=500e-9 W=3e-6
.ends SAVM1427

.subckt SAVM1428 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3028 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1428 L=500e-9 W=3e-6
.ends SAVM1428

.subckt SAVM1429 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3029 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1429 L=500e-9 W=3e-6
.ends SAVM1429

.subckt SAVM1430 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3030 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1430 L=500e-9 W=3e-6
.ends SAVM1430

.subckt SAVM1431 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3031 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1431 L=500e-9 W=3e-6
.ends SAVM1431

.subckt SAVM1432 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3032 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1432 L=500e-9 W=3e-6
.ends SAVM1432

.subckt SAVM1433 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3033 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1433 L=500e-9 W=3e-6
.ends SAVM1433

.subckt SAVM1434 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3034 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1434 L=500e-9 W=3e-6
.ends SAVM1434

.subckt SAVM1435 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3035 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1435 L=500e-9 W=3e-6
.ends SAVM1435

.subckt SAVM1436 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3036 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1436 L=500e-9 W=3e-6
.ends SAVM1436

.subckt SAVM1437 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3037 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1437 L=500e-9 W=3e-6
.ends SAVM1437

.subckt SAVM1438 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3038 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1438 L=500e-9 W=3e-6
.ends SAVM1438

.subckt SAVM1439 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3039 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1439 L=500e-9 W=3e-6
.ends SAVM1439

.subckt SAVM1440 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3040 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1440 L=500e-9 W=3e-6
.ends SAVM1440

.subckt SAVM1441 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3041 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1441 L=500e-9 W=3e-6
.ends SAVM1441

.subckt SAVM1442 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3042 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1442 L=500e-9 W=3e-6
.ends SAVM1442

.subckt SAVM1443 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3043 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1443 L=500e-9 W=3e-6
.ends SAVM1443

.subckt SAVM1444 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3044 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1444 L=500e-9 W=3e-6
.ends SAVM1444

.subckt SAVM1445 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3045 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1445 L=500e-9 W=3e-6
.ends SAVM1445

.subckt SAVM1446 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3046 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1446 L=500e-9 W=3e-6
.ends SAVM1446

.subckt SAVM1447 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3047 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1447 L=500e-9 W=3e-6
.ends SAVM1447

.subckt SAVM1448 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3048 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1448 L=500e-9 W=3e-6
.ends SAVM1448

.subckt SAVM1449 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3049 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1449 L=500e-9 W=3e-6
.ends SAVM1449

.subckt SAVM1450 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3050 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1450 L=500e-9 W=3e-6
.ends SAVM1450

.subckt SAVM1451 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3051 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1451 L=500e-9 W=3e-6
.ends SAVM1451

.subckt SAVM1452 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3052 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1452 L=500e-9 W=3e-6
.ends SAVM1452

.subckt SAVM1453 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3053 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1453 L=500e-9 W=3e-6
.ends SAVM1453

.subckt SAVM1454 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3054 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1454 L=500e-9 W=3e-6
.ends SAVM1454

.subckt SAVM1455 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3055 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1455 L=500e-9 W=3e-6
.ends SAVM1455

.subckt SAVM1456 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3056 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1456 L=500e-9 W=3e-6
.ends SAVM1456

.subckt SAVM1457 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3057 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1457 L=500e-9 W=3e-6
.ends SAVM1457

.subckt SAVM1458 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3058 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1458 L=500e-9 W=3e-6
.ends SAVM1458

.subckt SAVM1459 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3059 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1459 L=500e-9 W=3e-6
.ends SAVM1459

.subckt SAVM1460 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3060 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1460 L=500e-9 W=3e-6
.ends SAVM1460

.subckt SAVM1461 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3061 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1461 L=500e-9 W=3e-6
.ends SAVM1461

.subckt SAVM1462 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3062 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1462 L=500e-9 W=3e-6
.ends SAVM1462

.subckt SAVM1463 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3063 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1463 L=500e-9 W=3e-6
.ends SAVM1463

.subckt SAVM1464 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3064 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1464 L=500e-9 W=3e-6
.ends SAVM1464

.subckt SAVM1465 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3065 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1465 L=500e-9 W=3e-6
.ends SAVM1465

.subckt SAVM1466 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3066 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1466 L=500e-9 W=3e-6
.ends SAVM1466

.subckt SAVM1467 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3067 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1467 L=500e-9 W=3e-6
.ends SAVM1467

.subckt SAVM1468 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3068 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1468 L=500e-9 W=3e-6
.ends SAVM1468

.subckt SAVM1469 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3069 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1469 L=500e-9 W=3e-6
.ends SAVM1469

.subckt SAVM1470 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3070 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1470 L=500e-9 W=3e-6
.ends SAVM1470

.subckt SAVM1471 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3071 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1471 L=500e-9 W=3e-6
.ends SAVM1471

.subckt SAVM1472 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3072 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1472 L=500e-9 W=3e-6
.ends SAVM1472

.subckt SAVM1473 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3073 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1473 L=500e-9 W=3e-6
.ends SAVM1473

.subckt SAVM1474 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3074 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1474 L=500e-9 W=3e-6
.ends SAVM1474

.subckt SAVM1475 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3075 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1475 L=500e-9 W=3e-6
.ends SAVM1475

.subckt SAVM1476 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3076 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1476 L=500e-9 W=3e-6
.ends SAVM1476

.subckt SAVM1477 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3077 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1477 L=500e-9 W=3e-6
.ends SAVM1477

.subckt SAVM1478 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3078 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1478 L=500e-9 W=3e-6
.ends SAVM1478

.subckt SAVM1479 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3079 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1479 L=500e-9 W=3e-6
.ends SAVM1479

.subckt SAVM1480 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3080 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1480 L=500e-9 W=3e-6
.ends SAVM1480

.subckt SAVM1481 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3081 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1481 L=500e-9 W=3e-6
.ends SAVM1481

.subckt SAVM1482 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3082 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1482 L=500e-9 W=3e-6
.ends SAVM1482

.subckt SAVM1483 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3083 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1483 L=500e-9 W=3e-6
.ends SAVM1483

.subckt SAVM1484 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3084 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1484 L=500e-9 W=3e-6
.ends SAVM1484

.subckt SAVM1485 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3085 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1485 L=500e-9 W=3e-6
.ends SAVM1485

.subckt SAVM1486 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3086 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1486 L=500e-9 W=3e-6
.ends SAVM1486

.subckt SAVM1487 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3087 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1487 L=500e-9 W=3e-6
.ends SAVM1487

.subckt SAVM1488 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3088 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1488 L=500e-9 W=3e-6
.ends SAVM1488

.subckt SAVM1489 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3089 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1489 L=500e-9 W=3e-6
.ends SAVM1489

.subckt SAVM1490 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3090 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1490 L=500e-9 W=3e-6
.ends SAVM1490

.subckt SAVM1491 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3091 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1491 L=500e-9 W=3e-6
.ends SAVM1491

.subckt SAVM1492 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3092 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1492 L=500e-9 W=3e-6
.ends SAVM1492

.subckt SAVM1493 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3093 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1493 L=500e-9 W=3e-6
.ends SAVM1493

.subckt SAVM1494 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3094 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1494 L=500e-9 W=3e-6
.ends SAVM1494

.subckt SAVM1495 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3095 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1495 L=500e-9 W=3e-6
.ends SAVM1495

.subckt SAVM1496 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3096 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1496 L=500e-9 W=3e-6
.ends SAVM1496

.subckt SAVM1497 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3097 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1497 L=500e-9 W=3e-6
.ends SAVM1497

.subckt SAVM1498 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3098 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1498 L=500e-9 W=3e-6
.ends SAVM1498

.subckt SAVM1499 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3099 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1499 L=500e-9 W=3e-6
.ends SAVM1499

.subckt SAVM1500 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3100 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1500 L=500e-9 W=3e-6
.ends SAVM1500

.subckt SAVM1501 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3101 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1501 L=500e-9 W=3e-6
.ends SAVM1501

.subckt SAVM1502 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3102 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1502 L=500e-9 W=3e-6
.ends SAVM1502

.subckt SAVM1503 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3103 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1503 L=500e-9 W=3e-6
.ends SAVM1503

.subckt SAVM1504 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3104 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1504 L=500e-9 W=3e-6
.ends SAVM1504

.subckt SAVM1505 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3105 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1505 L=500e-9 W=3e-6
.ends SAVM1505

.subckt SAVM1506 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3106 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1506 L=500e-9 W=3e-6
.ends SAVM1506

.subckt SAVM1507 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3107 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1507 L=500e-9 W=3e-6
.ends SAVM1507

.subckt SAVM1508 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3108 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1508 L=500e-9 W=3e-6
.ends SAVM1508

.subckt SAVM1509 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3109 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1509 L=500e-9 W=3e-6
.ends SAVM1509

.subckt SAVM1510 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3110 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1510 L=500e-9 W=3e-6
.ends SAVM1510

.subckt SAVM1511 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3111 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1511 L=500e-9 W=3e-6
.ends SAVM1511

.subckt SAVM1512 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3112 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1512 L=500e-9 W=3e-6
.ends SAVM1512

.subckt SAVM1513 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3113 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1513 L=500e-9 W=3e-6
.ends SAVM1513

.subckt SAVM1514 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3114 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1514 L=500e-9 W=3e-6
.ends SAVM1514

.subckt SAVM1515 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3115 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1515 L=500e-9 W=3e-6
.ends SAVM1515

.subckt SAVM1516 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3116 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1516 L=500e-9 W=3e-6
.ends SAVM1516

.subckt SAVM1517 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3117 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1517 L=500e-9 W=3e-6
.ends SAVM1517

.subckt SAVM1518 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3118 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1518 L=500e-9 W=3e-6
.ends SAVM1518

.subckt SAVM1519 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3119 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1519 L=500e-9 W=3e-6
.ends SAVM1519

.subckt SAVM1520 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3120 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1520 L=500e-9 W=3e-6
.ends SAVM1520

.subckt SAVM1521 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3121 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1521 L=500e-9 W=3e-6
.ends SAVM1521

.subckt SAVM1522 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3122 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1522 L=500e-9 W=3e-6
.ends SAVM1522

.subckt SAVM1523 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3123 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1523 L=500e-9 W=3e-6
.ends SAVM1523

.subckt SAVM1524 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3124 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1524 L=500e-9 W=3e-6
.ends SAVM1524

.subckt SAVM1525 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3125 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1525 L=500e-9 W=3e-6
.ends SAVM1525

.subckt SAVM1526 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3126 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1526 L=500e-9 W=3e-6
.ends SAVM1526

.subckt SAVM1527 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3127 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1527 L=500e-9 W=3e-6
.ends SAVM1527

.subckt SAVM1528 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3128 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1528 L=500e-9 W=3e-6
.ends SAVM1528

.subckt SAVM1529 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3129 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1529 L=500e-9 W=3e-6
.ends SAVM1529

.subckt SAVM1530 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3130 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1530 L=500e-9 W=3e-6
.ends SAVM1530

.subckt SAVM1531 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3131 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1531 L=500e-9 W=3e-6
.ends SAVM1531

.subckt SAVM1532 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3132 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1532 L=500e-9 W=3e-6
.ends SAVM1532

.subckt SAVM1533 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3133 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1533 L=500e-9 W=3e-6
.ends SAVM1533

.subckt SAVM1534 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3134 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1534 L=500e-9 W=3e-6
.ends SAVM1534

.subckt SAVM1535 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3135 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1535 L=500e-9 W=3e-6
.ends SAVM1535

.subckt SAVM1536 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3136 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1536 L=500e-9 W=3e-6
.ends SAVM1536

.subckt SAVM1537 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3137 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1537 L=500e-9 W=3e-6
.ends SAVM1537

.subckt SAVM1538 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3138 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1538 L=500e-9 W=3e-6
.ends SAVM1538

.subckt SAVM1539 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3139 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1539 L=500e-9 W=3e-6
.ends SAVM1539

.subckt SAVM1540 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3140 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1540 L=500e-9 W=3e-6
.ends SAVM1540

.subckt SAVM1541 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3141 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1541 L=500e-9 W=3e-6
.ends SAVM1541

.subckt SAVM1542 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3142 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1542 L=500e-9 W=3e-6
.ends SAVM1542

.subckt SAVM1543 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3143 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1543 L=500e-9 W=3e-6
.ends SAVM1543

.subckt SAVM1544 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3144 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1544 L=500e-9 W=3e-6
.ends SAVM1544

.subckt SAVM1545 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3145 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1545 L=500e-9 W=3e-6
.ends SAVM1545

.subckt SAVM1546 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3146 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1546 L=500e-9 W=3e-6
.ends SAVM1546

.subckt SAVM1547 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3147 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1547 L=500e-9 W=3e-6
.ends SAVM1547

.subckt SAVM1548 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3148 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1548 L=500e-9 W=3e-6
.ends SAVM1548

.subckt SAVM1549 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3149 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1549 L=500e-9 W=3e-6
.ends SAVM1549

.subckt SAVM1550 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3150 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1550 L=500e-9 W=3e-6
.ends SAVM1550

.subckt SAVM1551 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3151 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1551 L=500e-9 W=3e-6
.ends SAVM1551

.subckt SAVM1552 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3152 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1552 L=500e-9 W=3e-6
.ends SAVM1552

.subckt SAVM1553 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3153 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1553 L=500e-9 W=3e-6
.ends SAVM1553

.subckt SAVM1554 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3154 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1554 L=500e-9 W=3e-6
.ends SAVM1554

.subckt SAVM1555 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3155 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1555 L=500e-9 W=3e-6
.ends SAVM1555

.subckt SAVM1556 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3156 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1556 L=500e-9 W=3e-6
.ends SAVM1556

.subckt SAVM1557 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3157 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1557 L=500e-9 W=3e-6
.ends SAVM1557

.subckt SAVM1558 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3158 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1558 L=500e-9 W=3e-6
.ends SAVM1558

.subckt SAVM1559 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3159 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1559 L=500e-9 W=3e-6
.ends SAVM1559

.subckt SAVM1560 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3160 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1560 L=500e-9 W=3e-6
.ends SAVM1560

.subckt SAVM1561 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3161 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1561 L=500e-9 W=3e-6
.ends SAVM1561

.subckt SAVM1562 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3162 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1562 L=500e-9 W=3e-6
.ends SAVM1562

.subckt SAVM1563 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3163 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1563 L=500e-9 W=3e-6
.ends SAVM1563

.subckt SAVM1564 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3164 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1564 L=500e-9 W=3e-6
.ends SAVM1564

.subckt SAVM1565 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3165 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1565 L=500e-9 W=3e-6
.ends SAVM1565

.subckt SAVM1566 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3166 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1566 L=500e-9 W=3e-6
.ends SAVM1566

.subckt SAVM1567 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3167 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1567 L=500e-9 W=3e-6
.ends SAVM1567

.subckt SAVM1568 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3168 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1568 L=500e-9 W=3e-6
.ends SAVM1568

.subckt SAVM1569 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3169 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1569 L=500e-9 W=3e-6
.ends SAVM1569

.subckt SAVM1570 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3170 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1570 L=500e-9 W=3e-6
.ends SAVM1570

.subckt SAVM1571 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3171 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1571 L=500e-9 W=3e-6
.ends SAVM1571

.subckt SAVM1572 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3172 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1572 L=500e-9 W=3e-6
.ends SAVM1572

.subckt SAVM1573 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3173 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1573 L=500e-9 W=3e-6
.ends SAVM1573

.subckt SAVM1574 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3174 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1574 L=500e-9 W=3e-6
.ends SAVM1574

.subckt SAVM1575 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3175 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1575 L=500e-9 W=3e-6
.ends SAVM1575

.subckt SAVM1576 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3176 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1576 L=500e-9 W=3e-6
.ends SAVM1576

.subckt SAVM1577 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3177 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1577 L=500e-9 W=3e-6
.ends SAVM1577

.subckt SAVM1578 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3178 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1578 L=500e-9 W=3e-6
.ends SAVM1578

.subckt SAVM1579 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3179 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1579 L=500e-9 W=3e-6
.ends SAVM1579

.subckt SAVM1580 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3180 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1580 L=500e-9 W=3e-6
.ends SAVM1580

.subckt SAVM1581 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3181 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1581 L=500e-9 W=3e-6
.ends SAVM1581

.subckt SAVM1582 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3182 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1582 L=500e-9 W=3e-6
.ends SAVM1582

.subckt SAVM1583 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3183 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1583 L=500e-9 W=3e-6
.ends SAVM1583

.subckt SAVM1584 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3184 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1584 L=500e-9 W=3e-6
.ends SAVM1584

.subckt SAVM1585 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3185 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1585 L=500e-9 W=3e-6
.ends SAVM1585

.subckt SAVM1586 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3186 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1586 L=500e-9 W=3e-6
.ends SAVM1586

.subckt SAVM1587 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3187 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1587 L=500e-9 W=3e-6
.ends SAVM1587

.subckt SAVM1588 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3188 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1588 L=500e-9 W=3e-6
.ends SAVM1588

.subckt SAVM1589 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3189 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1589 L=500e-9 W=3e-6
.ends SAVM1589

.subckt SAVM1590 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3190 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1590 L=500e-9 W=3e-6
.ends SAVM1590

.subckt SAVM1591 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3191 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1591 L=500e-9 W=3e-6
.ends SAVM1591

.subckt SAVM1592 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3192 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1592 L=500e-9 W=3e-6
.ends SAVM1592

.subckt SAVM1593 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3193 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1593 L=500e-9 W=3e-6
.ends SAVM1593

.subckt SAVM1594 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3194 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1594 L=500e-9 W=3e-6
.ends SAVM1594

.subckt SAVM1595 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3195 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1595 L=500e-9 W=3e-6
.ends SAVM1595

.subckt SAVM1596 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3196 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1596 L=500e-9 W=3e-6
.ends SAVM1596

.subckt SAVM1597 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3197 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1597 L=500e-9 W=3e-6
.ends SAVM1597

.subckt SAVM1598 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3198 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1598 L=500e-9 W=3e-6
.ends SAVM1598

.subckt SAVM1599 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3199 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1599 L=500e-9 W=3e-6
.ends SAVM1599

.subckt SAVM1600 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3200 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1600 L=500e-9 W=3e-6
.ends SAVM1600

.subckt SAVM1601 bl blb dl vdd
m1 dl net19 vdd vdd P L=180e-9 W=1e-6
m0 net19 net19 vdd vdd P L=180e-9 W=1e-6
m3 dl blb 0 0 N3201 L=500e-9 W=3e-6
m2 net19 bl 0 0 N1601 L=500e-9 W=3e-6
.ends SAVM1601

xl0b0c0 l0bl0 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b0c1 l0bl0 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b0c2 l0bl0 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b0c3 l0bl0 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b0c4 l0bl0 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b0c5 l0bl0 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b0c6 l0bl0 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b0c7 l0bl0 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b0c8 l0bl0 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b0c9 l0bl0 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b0c10 l0bl0 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b0c11 l0bl0 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b0c12 l0bl0 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b0c13 l0bl0 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b0c14 l0bl0 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b0c15 l0bl0 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b0c16 l0bl0 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b0c17 l0bl0 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b0c18 l0bl0 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b0c19 l0bl0 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b0c20 l0bl0 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b0c21 l0bl0 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b0c22 l0bl0 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b0c23 l0bl0 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b0c24 l0bl0 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b0c25 l0bl0 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b0c26 l0bl0 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b0c27 l0bl0 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b0c28 l0bl0 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b0c29 l0bl0 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b0c30 l0bl0 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b0c31 l0bl0 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b0c32 l0bl0 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b0c33 l0bl0 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b0c34 l0bl0 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b0c35 l0bl0 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b0c36 l0bl0 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b0c37 l0bl0 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b0c38 l0bl0 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b0c39 l0bl0 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b0c40 l0bl0 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b0c41 l0bl0 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b0c42 l0bl0 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b0c43 l0bl0 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b0c44 l0bl0 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b0c45 l0bl0 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b0c46 l0bl0 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b0c47 l0bl0 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b0c48 l0bl0 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b0c49 l0bl0 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b0c50 l0bl0 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b0c51 l0bl0 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b0c52 l0bl0 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b0c53 l0bl0 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b0c54 l0bl0 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b0c55 l0bl0 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b0c56 l0bl0 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b0c57 l0bl0 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b0c58 l0bl0 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b0c59 l0bl0 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b0c60 l0bl0 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b0c61 l0bl0 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b0c62 l0bl0 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b0c63 l0bl0 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b0c64 l0bl0 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b0c65 l0bl0 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b0c66 l0bl0 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b0c67 l0bl0 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b0c68 l0bl0 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b0c69 l0bl0 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b0c70 l0bl0 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b0c71 l0bl0 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b0c72 l0bl0 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b0c73 l0bl0 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b0c74 l0bl0 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b0c75 l0bl0 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b0c76 l0bl0 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b0c77 l0bl0 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b0c78 l0bl0 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b0c79 l0bl0 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b0c80 l0bl0 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b0c81 l0bl0 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b0c82 l0bl0 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b0c83 l0bl0 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b0c84 l0bl0 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b0c85 l0bl0 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b0c86 l0bl0 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b0c87 l0bl0 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b0c88 l0bl0 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b0c89 l0bl0 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b0c90 l0bl0 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b0c91 l0bl0 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b0c92 l0bl0 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b0c93 l0bl0 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b0c94 l0bl0 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b0c95 l0bl0 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b0c96 l0bl0 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b0c97 l0bl0 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b0c98 l0bl0 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b0c99 l0bl0 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b0c100 l0bl0 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b0c101 l0bl0 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b0c102 l0bl0 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b0c103 l0bl0 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b0c104 l0bl0 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b0c105 l0bl0 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b0c106 l0bl0 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b0c107 l0bl0 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b0c108 l0bl0 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b0c109 l0bl0 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b0c110 l0bl0 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b0c111 l0bl0 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b0c112 l0bl0 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b0c113 l0bl0 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b0c114 l0bl0 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b0c115 l0bl0 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b0c116 l0bl0 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b0c117 l0bl0 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b0c118 l0bl0 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b0c119 l0bl0 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b0c120 l0bl0 vdd x120 x120b CELLD r1=900e3 r0=10000e3
xl0b0c121 l0bl0 vdd x121 x121b CELLD r1=900e3 r0=10000e3
xl0b0c122 l0bl0 vdd x122 x122b CELLD r1=900e3 r0=10000e3
xl0b0c123 l0bl0 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b0c124 l0bl0 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b0c125 l0bl0 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b0c126 l0bl0 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b0c127 l0bl0 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b0c128 l0bl0 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b0c129 l0bl0 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b0c130 l0bl0 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b0c131 l0bl0 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b0c132 l0bl0 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b0c133 l0bl0 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b0c134 l0bl0 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b0c135 l0bl0 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b0c136 l0bl0 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b0c137 l0bl0 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b0c138 l0bl0 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b0c139 l0bl0 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b0c140 l0bl0 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b0c141 l0bl0 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b0c142 l0bl0 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b0c143 l0bl0 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b0c144 l0bl0 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b0c145 l0bl0 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b0c146 l0bl0 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b0c147 l0bl0 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b0c148 l0bl0 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b0c149 l0bl0 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b0c150 l0bl0 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b0c151 l0bl0 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b0c152 l0bl0 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b0c153 l0bl0 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b0c154 l0bl0 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b0c155 l0bl0 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b0c156 l0bl0 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b0c157 l0bl0 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b0c158 l0bl0 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b0c159 l0bl0 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b0c160 l0bl0 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b0c161 l0bl0 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b0c162 l0bl0 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b0c163 l0bl0 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b0c164 l0bl0 vdd x164 x164b CELLD r1=10000e3 r0=900e3
xl0b0c165 l0bl0 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b0c166 l0bl0 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b0c167 l0bl0 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b0c168 l0bl0 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b0c169 l0bl0 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b0c170 l0bl0 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b0c171 l0bl0 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b0c172 l0bl0 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b0c173 l0bl0 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b0c174 l0bl0 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b0c175 l0bl0 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b0c176 l0bl0 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b0c177 l0bl0 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b0c178 l0bl0 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b0c179 l0bl0 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b0c180 l0bl0 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b0c181 l0bl0 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b0c182 l0bl0 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b0c183 l0bl0 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b0c184 l0bl0 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b0c185 l0bl0 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b0c186 l0bl0 vdd x186 x186b CELLD r1=10000e3 r0=900e3
xl0b0c187 l0bl0 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b0c188 l0bl0 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b0c189 l0bl0 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b0c190 l0bl0 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b0c191 l0bl0 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b0c192 l0bl0 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b0c193 l0bl0 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b0c194 l0bl0 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b0c195 l0bl0 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b0c196 l0bl0 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b0c197 l0bl0 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b0c198 l0bl0 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b0c199 l0bl0 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b0c200 l0bl0 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b0c201 l0bl0 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b0c202 l0bl0 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b0c203 l0bl0 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b0c204 l0bl0 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b0c205 l0bl0 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b0c206 l0bl0 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b0c207 l0bl0 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b0c208 l0bl0 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b0c209 l0bl0 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b0c210 l0bl0 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b0c211 l0bl0 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b0c212 l0bl0 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b0c213 l0bl0 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b0c214 l0bl0 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b0c215 l0bl0 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b0c216 l0bl0 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b0c217 l0bl0 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b0c218 l0bl0 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b0c219 l0bl0 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b0c220 l0bl0 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b0c221 l0bl0 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b0c222 l0bl0 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b0c223 l0bl0 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b0c224 l0bl0 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b0c225 l0bl0 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b0c226 l0bl0 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b0c227 l0bl0 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b0c228 l0bl0 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b0c229 l0bl0 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b0c230 l0bl0 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b0c231 l0bl0 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b0c232 l0bl0 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b0c233 l0bl0 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b0c234 l0bl0 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b0c235 l0bl0 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b0c236 l0bl0 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b0c237 l0bl0 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b0c238 l0bl0 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b0c239 l0bl0 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b0c240 l0bl0 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b0c241 l0bl0 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b0c242 l0bl0 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b0c243 l0bl0 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b0c244 l0bl0 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b0c245 l0bl0 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b0c246 l0bl0 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b0c247 l0bl0 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b0c248 l0bl0 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b0c249 l0bl0 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b0c250 l0bl0 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b0c251 l0bl0 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b0c252 l0bl0 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b0c253 l0bl0 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b0c254 l0bl0 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b0c255 l0bl0 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b0c256 l0bl0 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b0c257 l0bl0 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b0c258 l0bl0 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b0c259 l0bl0 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b0c260 l0bl0 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b0c261 l0bl0 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b0c262 l0bl0 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b0c263 l0bl0 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b0c264 l0bl0 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b0c265 l0bl0 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b0c266 l0bl0 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b0c267 l0bl0 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b0c268 l0bl0 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b0c269 l0bl0 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b0c270 l0bl0 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b0c271 l0bl0 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b0c272 l0bl0 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b0c273 l0bl0 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b0c274 l0bl0 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b0c275 l0bl0 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b0c276 l0bl0 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b0c277 l0bl0 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b0c278 l0bl0 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b0c279 l0bl0 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b0c280 l0bl0 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b0c281 l0bl0 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b0c282 l0bl0 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b0c283 l0bl0 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b0c284 l0bl0 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b0c285 l0bl0 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b0c286 l0bl0 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b0c287 l0bl0 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b0c288 l0bl0 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b0c289 l0bl0 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b0c290 l0bl0 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b0c291 l0bl0 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b0c292 l0bl0 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b0c293 l0bl0 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b0c294 l0bl0 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b0c295 l0bl0 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b0c296 l0bl0 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b0c297 l0bl0 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b0c298 l0bl0 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b0c299 l0bl0 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b0c300 l0bl0 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b0c301 l0bl0 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b0c302 l0bl0 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b0c303 l0bl0 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b0c304 l0bl0 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b0c305 l0bl0 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b0c306 l0bl0 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b0c307 l0bl0 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b0c308 l0bl0 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b0c309 l0bl0 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b0c310 l0bl0 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b0c311 l0bl0 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b0c312 l0bl0 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b0c313 l0bl0 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b0c314 l0bl0 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b0c315 l0bl0 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b0c316 l0bl0 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b0c317 l0bl0 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b0c318 l0bl0 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b0c319 l0bl0 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b0c320 l0bl0 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b0c321 l0bl0 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b0c322 l0bl0 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b0c323 l0bl0 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b0c324 l0bl0 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b0c325 l0bl0 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b0c326 l0bl0 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b0c327 l0bl0 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b0c328 l0bl0 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b0c329 l0bl0 vdd x329 x329b CELLD r1=900e3 r0=10000e3
xl0b0c330 l0bl0 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b0c331 l0bl0 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b0c332 l0bl0 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b0c333 l0bl0 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b0c334 l0bl0 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b0c335 l0bl0 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b0c336 l0bl0 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b0c337 l0bl0 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b0c338 l0bl0 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b0c339 l0bl0 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b0c340 l0bl0 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b0c341 l0bl0 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b0c342 l0bl0 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b0c343 l0bl0 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b0c344 l0bl0 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b0c345 l0bl0 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b0c346 l0bl0 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b0c347 l0bl0 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b0c348 l0bl0 vdd x348 x348b CELLD r1=10000e3 r0=900e3
xl0b0c349 l0bl0 vdd x349 x349b CELLD r1=10000e3 r0=900e3
xl0b0c350 l0bl0 vdd x350 x350b CELLD r1=10000e3 r0=900e3
xl0b0c351 l0bl0 vdd x351 x351b CELLD r1=10000e3 r0=900e3
xl0b0c352 l0bl0 vdd x352 x352b CELLD r1=10000e3 r0=900e3
xl0b0c353 l0bl0 vdd x353 x353b CELLD r1=10000e3 r0=900e3
xl0b0c354 l0bl0 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b0c355 l0bl0 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b0c356 l0bl0 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b0c357 l0bl0 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b0c358 l0bl0 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b0c359 l0bl0 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b0c360 l0bl0 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b0c361 l0bl0 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b0c362 l0bl0 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b0c363 l0bl0 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b0c364 l0bl0 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b0c365 l0bl0 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b0c366 l0bl0 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b0c367 l0bl0 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b0c368 l0bl0 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b0c369 l0bl0 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b0c370 l0bl0 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b0c371 l0bl0 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b0c372 l0bl0 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b0c373 l0bl0 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b0c374 l0bl0 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b0c375 l0bl0 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b0c376 l0bl0 vdd x376 x376b CELLD r1=10000e3 r0=900e3
xl0b0c377 l0bl0 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b0c378 l0bl0 vdd x378 x378b CELLD r1=10000e3 r0=900e3
xl0b0c379 l0bl0 vdd x379 x379b CELLD r1=10000e3 r0=900e3
xl0b0c380 l0bl0 vdd x380 x380b CELLD r1=10000e3 r0=900e3
xl0b0c381 l0bl0 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b0c382 l0bl0 vdd x382 x382b CELLD r1=10000e3 r0=900e3
xl0b0c383 l0bl0 vdd x383 x383b CELLD r1=10000e3 r0=900e3
xl0b0c384 l0bl0 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b0c385 l0bl0 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b0c386 l0bl0 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b0c387 l0bl0 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b0c388 l0bl0 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b0c389 l0bl0 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b0c390 l0bl0 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b0c391 l0bl0 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b0c392 l0bl0 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b0c393 l0bl0 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b0c394 l0bl0 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b0c395 l0bl0 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b0c396 l0bl0 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b0c397 l0bl0 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b0c398 l0bl0 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b0c399 l0bl0 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b0c400 l0bl0 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b0c401 l0bl0 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b0c402 l0bl0 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b0c403 l0bl0 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b0c404 l0bl0 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b0c405 l0bl0 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b0c406 l0bl0 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b0c407 l0bl0 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b0c408 l0bl0 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b0c409 l0bl0 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b0c410 l0bl0 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b0c411 l0bl0 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b0c412 l0bl0 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b0c413 l0bl0 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b0c414 l0bl0 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b0c415 l0bl0 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b0c416 l0bl0 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b0c417 l0bl0 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b0c418 l0bl0 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b0c419 l0bl0 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b0c420 l0bl0 vdd x420 x420b CELLD r1=10000e3 r0=900e3
xl0b0c421 l0bl0 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b0c422 l0bl0 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b0c423 l0bl0 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b0c424 l0bl0 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b0c425 l0bl0 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b0c426 l0bl0 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b0c427 l0bl0 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b0c428 l0bl0 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b0c429 l0bl0 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b0c430 l0bl0 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b0c431 l0bl0 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b0c432 l0bl0 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b0c433 l0bl0 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b0c434 l0bl0 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b0c435 l0bl0 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b0c436 l0bl0 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b0c437 l0bl0 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b0c438 l0bl0 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b0c439 l0bl0 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b0c440 l0bl0 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b0c441 l0bl0 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b0c442 l0bl0 vdd x442 x442b CELLD r1=900e3 r0=10000e3
xl0b0c443 l0bl0 vdd x443 x443b CELLD r1=900e3 r0=10000e3
xl0b0c444 l0bl0 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b0c445 l0bl0 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b0c446 l0bl0 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b0c447 l0bl0 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b0c448 l0bl0 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b0c449 l0bl0 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b0c450 l0bl0 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b0c451 l0bl0 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b0c452 l0bl0 vdd x452 x452b CELLD r1=900e3 r0=10000e3
xl0b0c453 l0bl0 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b0c454 l0bl0 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b0c455 l0bl0 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b0c456 l0bl0 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b0c457 l0bl0 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b0c458 l0bl0 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b0c459 l0bl0 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b0c460 l0bl0 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b0c461 l0bl0 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b0c462 l0bl0 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b0c463 l0bl0 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b0c464 l0bl0 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b0c465 l0bl0 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b0c466 l0bl0 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b0c467 l0bl0 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b0c468 l0bl0 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b0c469 l0bl0 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b0c470 l0bl0 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b0c471 l0bl0 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b0c472 l0bl0 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b0c473 l0bl0 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b0c474 l0bl0 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b0c475 l0bl0 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b0c476 l0bl0 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b0c477 l0bl0 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b0c478 l0bl0 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b0c479 l0bl0 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b0c480 l0bl0 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b0c481 l0bl0 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b0c482 l0bl0 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b0c483 l0bl0 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b0c484 l0bl0 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b0c485 l0bl0 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b0c486 l0bl0 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b0c487 l0bl0 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b0c488 l0bl0 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b0c489 l0bl0 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b0c490 l0bl0 vdd x490 x490b CELLD r1=10000e3 r0=900e3
xl0b0c491 l0bl0 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b0c492 l0bl0 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b0c493 l0bl0 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b0c494 l0bl0 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b0c495 l0bl0 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b0c496 l0bl0 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b0c497 l0bl0 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b0c498 l0bl0 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b0c499 l0bl0 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b0c500 l0bl0 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b0c501 l0bl0 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b0c502 l0bl0 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b0c503 l0bl0 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b0c504 l0bl0 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b0c505 l0bl0 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b0c506 l0bl0 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b0c507 l0bl0 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b0c508 l0bl0 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b0c509 l0bl0 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b0c510 l0bl0 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b0c511 l0bl0 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b0c512 l0bl0 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b0c513 l0bl0 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b0c514 l0bl0 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b0c515 l0bl0 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b0c516 l0bl0 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b0c517 l0bl0 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b0c518 l0bl0 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b0c519 l0bl0 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b0c520 l0bl0 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b0c521 l0bl0 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b0c522 l0bl0 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b0c523 l0bl0 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b0c524 l0bl0 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b0c525 l0bl0 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b0c526 l0bl0 vdd x526 x526b CELLD r1=900e3 r0=10000e3
xl0b0c527 l0bl0 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b0c528 l0bl0 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b0c529 l0bl0 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b0c530 l0bl0 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b0c531 l0bl0 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b0c532 l0bl0 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b0c533 l0bl0 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b0c534 l0bl0 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b0c535 l0bl0 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b0c536 l0bl0 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b0c537 l0bl0 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b0c538 l0bl0 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b0c539 l0bl0 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b0c540 l0bl0 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b0c541 l0bl0 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b0c542 l0bl0 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b0c543 l0bl0 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b0c544 l0bl0 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b0c545 l0bl0 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b0c546 l0bl0 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b0c547 l0bl0 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b0c548 l0bl0 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b0c549 l0bl0 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b0c550 l0bl0 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b0c551 l0bl0 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b0c552 l0bl0 vdd x552 x552b CELLD r1=900e3 r0=10000e3
xl0b0c553 l0bl0 vdd x553 x553b CELLD r1=900e3 r0=10000e3
xl0b0c554 l0bl0 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b0c555 l0bl0 vdd x555 x555b CELLD r1=900e3 r0=10000e3
xl0b0c556 l0bl0 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b0c557 l0bl0 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b0c558 l0bl0 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b0c559 l0bl0 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b0c560 l0bl0 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b0c561 l0bl0 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b0c562 l0bl0 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b0c563 l0bl0 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b0c564 l0bl0 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b0c565 l0bl0 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b0c566 l0bl0 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b0c567 l0bl0 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b0c568 l0bl0 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b0c569 l0bl0 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b0c570 l0bl0 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b0c571 l0bl0 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b0c572 l0bl0 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b0c573 l0bl0 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b0c574 l0bl0 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b0c575 l0bl0 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b0c576 l0bl0 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b0c577 l0bl0 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b0c578 l0bl0 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b0c579 l0bl0 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b0c580 l0bl0 vdd x580 x580b CELLD r1=900e3 r0=10000e3
xl0b0c581 l0bl0 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b0c582 l0bl0 vdd x582 x582b CELLD r1=900e3 r0=10000e3
xl0b0c583 l0bl0 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b0c584 l0bl0 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b0c585 l0bl0 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b0c586 l0bl0 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b0c587 l0bl0 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b0c588 l0bl0 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b0c589 l0bl0 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b0c590 l0bl0 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b0c591 l0bl0 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b0c592 l0bl0 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b0c593 l0bl0 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b0c594 l0bl0 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b0c595 l0bl0 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b0c596 l0bl0 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b0c597 l0bl0 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b0c598 l0bl0 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b0c599 l0bl0 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b0c600 l0bl0 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b0c601 l0bl0 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b0c602 l0bl0 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b0c603 l0bl0 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b0c604 l0bl0 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b0c605 l0bl0 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b0c606 l0bl0 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b0c607 l0bl0 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b0c608 l0bl0 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b0c609 l0bl0 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b0c610 l0bl0 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b0c611 l0bl0 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b0c612 l0bl0 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b0c613 l0bl0 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b0c614 l0bl0 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b0c615 l0bl0 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b0c616 l0bl0 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b0c617 l0bl0 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b0c618 l0bl0 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b0c619 l0bl0 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b0c620 l0bl0 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b0c621 l0bl0 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b0c622 l0bl0 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b0c623 l0bl0 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b0c624 l0bl0 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b0c625 l0bl0 vdd x625 x625b CELLD r1=900e3 r0=10000e3
xl0b0c626 l0bl0 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b0c627 l0bl0 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b0c628 l0bl0 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b0c629 l0bl0 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b0c630 l0bl0 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b0c631 l0bl0 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b0c632 l0bl0 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b0c633 l0bl0 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b0c634 l0bl0 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b0c635 l0bl0 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b0c636 l0bl0 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b0c637 l0bl0 vdd x637 x637b CELLD r1=10000e3 r0=900e3
xl0b0c638 l0bl0 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b0c639 l0bl0 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b0c640 l0bl0 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b0c641 l0bl0 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b0c642 l0bl0 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b0c643 l0bl0 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b0c644 l0bl0 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b0c645 l0bl0 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b0c646 l0bl0 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b0c647 l0bl0 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b0c648 l0bl0 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b0c649 l0bl0 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b0c650 l0bl0 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b0c651 l0bl0 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b0c652 l0bl0 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b0c653 l0bl0 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b0c654 l0bl0 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b0c655 l0bl0 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b0c656 l0bl0 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b0c657 l0bl0 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b0c658 l0bl0 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b0c659 l0bl0 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b0c660 l0bl0 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b0c661 l0bl0 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b0c662 l0bl0 vdd x662 x662b CELLD r1=10000e3 r0=900e3
xl0b0c663 l0bl0 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b0c664 l0bl0 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b0c665 l0bl0 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b0c666 l0bl0 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b0c667 l0bl0 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b0c668 l0bl0 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b0c669 l0bl0 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b0c670 l0bl0 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b0c671 l0bl0 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b0c672 l0bl0 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b0c673 l0bl0 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b0c674 l0bl0 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b0c675 l0bl0 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b0c676 l0bl0 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b0c677 l0bl0 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b0c678 l0bl0 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b0c679 l0bl0 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b0c680 l0bl0 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b0c681 l0bl0 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b0c682 l0bl0 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b0c683 l0bl0 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b0c684 l0bl0 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b0c685 l0bl0 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b0c686 l0bl0 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b0c687 l0bl0 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b0c688 l0bl0 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b0c689 l0bl0 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b0c690 l0bl0 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b0c691 l0bl0 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b0c692 l0bl0 vdd x692 x692b CELLD r1=10000e3 r0=900e3
xl0b0c693 l0bl0 vdd x693 x693b CELLD r1=10000e3 r0=900e3
xl0b0c694 l0bl0 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b0c695 l0bl0 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b0c696 l0bl0 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b0c697 l0bl0 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b0c698 l0bl0 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b0c699 l0bl0 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b0c700 l0bl0 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b0c701 l0bl0 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b0c702 l0bl0 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b0c703 l0bl0 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b0c704 l0bl0 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b0c705 l0bl0 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b0c706 l0bl0 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b0c707 l0bl0 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b0c708 l0bl0 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b0c709 l0bl0 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b0c710 l0bl0 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b0c711 l0bl0 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b0c712 l0bl0 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b0c713 l0bl0 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b0c714 l0bl0 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b0c715 l0bl0 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b0c716 l0bl0 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b0c717 l0bl0 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b0c718 l0bl0 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b0c719 l0bl0 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b0c720 l0bl0 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b0c721 l0bl0 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b0c722 l0bl0 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b0c723 l0bl0 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b0c724 l0bl0 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b0c725 l0bl0 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b0c726 l0bl0 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b0c727 l0bl0 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b0c728 l0bl0 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b0c729 l0bl0 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b0c730 l0bl0 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b0c731 l0bl0 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b0c732 l0bl0 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b0c733 l0bl0 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b0c734 l0bl0 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b0c735 l0bl0 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b0c736 l0bl0 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b0c737 l0bl0 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b0c738 l0bl0 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b0c739 l0bl0 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b0c740 l0bl0 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b0c741 l0bl0 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b0c742 l0bl0 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b0c743 l0bl0 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b0c744 l0bl0 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b0c745 l0bl0 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b0c746 l0bl0 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b0c747 l0bl0 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b0c748 l0bl0 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b0c749 l0bl0 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b0c750 l0bl0 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b0c751 l0bl0 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b0c752 l0bl0 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b0c753 l0bl0 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b0c754 l0bl0 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b0c755 l0bl0 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b0c756 l0bl0 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b0c757 l0bl0 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b0c758 l0bl0 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b0c759 l0bl0 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b0c760 l0bl0 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b0c761 l0bl0 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b0c762 l0bl0 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b0c763 l0bl0 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b0c764 l0bl0 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b0c765 l0bl0 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b0c766 l0bl0 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b0c767 l0bl0 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b0c768 l0bl0 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b0c769 l0bl0 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b0c770 l0bl0 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b0c771 l0bl0 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b0c772 l0bl0 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b0c773 l0bl0 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b0c774 l0bl0 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b0c775 l0bl0 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b0c776 l0bl0 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b0c777 l0bl0 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b0c778 l0bl0 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b0c779 l0bl0 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b0c780 l0bl0 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b0c781 l0bl0 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b0c782 l0bl0 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b0c783 l0bl0 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b1c0 l0bl1 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b1c1 l0bl1 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b1c2 l0bl1 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b1c3 l0bl1 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b1c4 l0bl1 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b1c5 l0bl1 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b1c6 l0bl1 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b1c7 l0bl1 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b1c8 l0bl1 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b1c9 l0bl1 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b1c10 l0bl1 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b1c11 l0bl1 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b1c12 l0bl1 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b1c13 l0bl1 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b1c14 l0bl1 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b1c15 l0bl1 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b1c16 l0bl1 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b1c17 l0bl1 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b1c18 l0bl1 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b1c19 l0bl1 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b1c20 l0bl1 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b1c21 l0bl1 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b1c22 l0bl1 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b1c23 l0bl1 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b1c24 l0bl1 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b1c25 l0bl1 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b1c26 l0bl1 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b1c27 l0bl1 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b1c28 l0bl1 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b1c29 l0bl1 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b1c30 l0bl1 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b1c31 l0bl1 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b1c32 l0bl1 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b1c33 l0bl1 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b1c34 l0bl1 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b1c35 l0bl1 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b1c36 l0bl1 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b1c37 l0bl1 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b1c38 l0bl1 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b1c39 l0bl1 vdd x39 x39b CELLD r1=10000e3 r0=900e3
xl0b1c40 l0bl1 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b1c41 l0bl1 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b1c42 l0bl1 vdd x42 x42b CELLD r1=10000e3 r0=900e3
xl0b1c43 l0bl1 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b1c44 l0bl1 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b1c45 l0bl1 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b1c46 l0bl1 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b1c47 l0bl1 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b1c48 l0bl1 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b1c49 l0bl1 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b1c50 l0bl1 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b1c51 l0bl1 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b1c52 l0bl1 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b1c53 l0bl1 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b1c54 l0bl1 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b1c55 l0bl1 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b1c56 l0bl1 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b1c57 l0bl1 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b1c58 l0bl1 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b1c59 l0bl1 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b1c60 l0bl1 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b1c61 l0bl1 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b1c62 l0bl1 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b1c63 l0bl1 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b1c64 l0bl1 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b1c65 l0bl1 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b1c66 l0bl1 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b1c67 l0bl1 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b1c68 l0bl1 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b1c69 l0bl1 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b1c70 l0bl1 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b1c71 l0bl1 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b1c72 l0bl1 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b1c73 l0bl1 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b1c74 l0bl1 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b1c75 l0bl1 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b1c76 l0bl1 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b1c77 l0bl1 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b1c78 l0bl1 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b1c79 l0bl1 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b1c80 l0bl1 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b1c81 l0bl1 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b1c82 l0bl1 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b1c83 l0bl1 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b1c84 l0bl1 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b1c85 l0bl1 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b1c86 l0bl1 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b1c87 l0bl1 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b1c88 l0bl1 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b1c89 l0bl1 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b1c90 l0bl1 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b1c91 l0bl1 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b1c92 l0bl1 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b1c93 l0bl1 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b1c94 l0bl1 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b1c95 l0bl1 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b1c96 l0bl1 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b1c97 l0bl1 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b1c98 l0bl1 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b1c99 l0bl1 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b1c100 l0bl1 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b1c101 l0bl1 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b1c102 l0bl1 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b1c103 l0bl1 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b1c104 l0bl1 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b1c105 l0bl1 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b1c106 l0bl1 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b1c107 l0bl1 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b1c108 l0bl1 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b1c109 l0bl1 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b1c110 l0bl1 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b1c111 l0bl1 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b1c112 l0bl1 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b1c113 l0bl1 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b1c114 l0bl1 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b1c115 l0bl1 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b1c116 l0bl1 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b1c117 l0bl1 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b1c118 l0bl1 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b1c119 l0bl1 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b1c120 l0bl1 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b1c121 l0bl1 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b1c122 l0bl1 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b1c123 l0bl1 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b1c124 l0bl1 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b1c125 l0bl1 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b1c126 l0bl1 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b1c127 l0bl1 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b1c128 l0bl1 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b1c129 l0bl1 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b1c130 l0bl1 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b1c131 l0bl1 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b1c132 l0bl1 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b1c133 l0bl1 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b1c134 l0bl1 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b1c135 l0bl1 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b1c136 l0bl1 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b1c137 l0bl1 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b1c138 l0bl1 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b1c139 l0bl1 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b1c140 l0bl1 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b1c141 l0bl1 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b1c142 l0bl1 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b1c143 l0bl1 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b1c144 l0bl1 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b1c145 l0bl1 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b1c146 l0bl1 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b1c147 l0bl1 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b1c148 l0bl1 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b1c149 l0bl1 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b1c150 l0bl1 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b1c151 l0bl1 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b1c152 l0bl1 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b1c153 l0bl1 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b1c154 l0bl1 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b1c155 l0bl1 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b1c156 l0bl1 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b1c157 l0bl1 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b1c158 l0bl1 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b1c159 l0bl1 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b1c160 l0bl1 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b1c161 l0bl1 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b1c162 l0bl1 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b1c163 l0bl1 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b1c164 l0bl1 vdd x164 x164b CELLD r1=10000e3 r0=900e3
xl0b1c165 l0bl1 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b1c166 l0bl1 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b1c167 l0bl1 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b1c168 l0bl1 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b1c169 l0bl1 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b1c170 l0bl1 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b1c171 l0bl1 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b1c172 l0bl1 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b1c173 l0bl1 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b1c174 l0bl1 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b1c175 l0bl1 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b1c176 l0bl1 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b1c177 l0bl1 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b1c178 l0bl1 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b1c179 l0bl1 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b1c180 l0bl1 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b1c181 l0bl1 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b1c182 l0bl1 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b1c183 l0bl1 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b1c184 l0bl1 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b1c185 l0bl1 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b1c186 l0bl1 vdd x186 x186b CELLD r1=10000e3 r0=900e3
xl0b1c187 l0bl1 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b1c188 l0bl1 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b1c189 l0bl1 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b1c190 l0bl1 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b1c191 l0bl1 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b1c192 l0bl1 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b1c193 l0bl1 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b1c194 l0bl1 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b1c195 l0bl1 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b1c196 l0bl1 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b1c197 l0bl1 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b1c198 l0bl1 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b1c199 l0bl1 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b1c200 l0bl1 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b1c201 l0bl1 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b1c202 l0bl1 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b1c203 l0bl1 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b1c204 l0bl1 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b1c205 l0bl1 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b1c206 l0bl1 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b1c207 l0bl1 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b1c208 l0bl1 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b1c209 l0bl1 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b1c210 l0bl1 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b1c211 l0bl1 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b1c212 l0bl1 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b1c213 l0bl1 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b1c214 l0bl1 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b1c215 l0bl1 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b1c216 l0bl1 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b1c217 l0bl1 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b1c218 l0bl1 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b1c219 l0bl1 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b1c220 l0bl1 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b1c221 l0bl1 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b1c222 l0bl1 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b1c223 l0bl1 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b1c224 l0bl1 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b1c225 l0bl1 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b1c226 l0bl1 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b1c227 l0bl1 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b1c228 l0bl1 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b1c229 l0bl1 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b1c230 l0bl1 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b1c231 l0bl1 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b1c232 l0bl1 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b1c233 l0bl1 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b1c234 l0bl1 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b1c235 l0bl1 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b1c236 l0bl1 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b1c237 l0bl1 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b1c238 l0bl1 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b1c239 l0bl1 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b1c240 l0bl1 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b1c241 l0bl1 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b1c242 l0bl1 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b1c243 l0bl1 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b1c244 l0bl1 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b1c245 l0bl1 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b1c246 l0bl1 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b1c247 l0bl1 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b1c248 l0bl1 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b1c249 l0bl1 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b1c250 l0bl1 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b1c251 l0bl1 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b1c252 l0bl1 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b1c253 l0bl1 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b1c254 l0bl1 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b1c255 l0bl1 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b1c256 l0bl1 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b1c257 l0bl1 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b1c258 l0bl1 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b1c259 l0bl1 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b1c260 l0bl1 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b1c261 l0bl1 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b1c262 l0bl1 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b1c263 l0bl1 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b1c264 l0bl1 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b1c265 l0bl1 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b1c266 l0bl1 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b1c267 l0bl1 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b1c268 l0bl1 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b1c269 l0bl1 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b1c270 l0bl1 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b1c271 l0bl1 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b1c272 l0bl1 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b1c273 l0bl1 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b1c274 l0bl1 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b1c275 l0bl1 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b1c276 l0bl1 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b1c277 l0bl1 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b1c278 l0bl1 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b1c279 l0bl1 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b1c280 l0bl1 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b1c281 l0bl1 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b1c282 l0bl1 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b1c283 l0bl1 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b1c284 l0bl1 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b1c285 l0bl1 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b1c286 l0bl1 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b1c287 l0bl1 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b1c288 l0bl1 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b1c289 l0bl1 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b1c290 l0bl1 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b1c291 l0bl1 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b1c292 l0bl1 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b1c293 l0bl1 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b1c294 l0bl1 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b1c295 l0bl1 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b1c296 l0bl1 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b1c297 l0bl1 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b1c298 l0bl1 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b1c299 l0bl1 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b1c300 l0bl1 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b1c301 l0bl1 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b1c302 l0bl1 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b1c303 l0bl1 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b1c304 l0bl1 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b1c305 l0bl1 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b1c306 l0bl1 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b1c307 l0bl1 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b1c308 l0bl1 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b1c309 l0bl1 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b1c310 l0bl1 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b1c311 l0bl1 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b1c312 l0bl1 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b1c313 l0bl1 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b1c314 l0bl1 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b1c315 l0bl1 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b1c316 l0bl1 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b1c317 l0bl1 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b1c318 l0bl1 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b1c319 l0bl1 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b1c320 l0bl1 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b1c321 l0bl1 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b1c322 l0bl1 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b1c323 l0bl1 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b1c324 l0bl1 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b1c325 l0bl1 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b1c326 l0bl1 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b1c327 l0bl1 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b1c328 l0bl1 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b1c329 l0bl1 vdd x329 x329b CELLD r1=900e3 r0=10000e3
xl0b1c330 l0bl1 vdd x330 x330b CELLD r1=900e3 r0=10000e3
xl0b1c331 l0bl1 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b1c332 l0bl1 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b1c333 l0bl1 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b1c334 l0bl1 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b1c335 l0bl1 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b1c336 l0bl1 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b1c337 l0bl1 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b1c338 l0bl1 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b1c339 l0bl1 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b1c340 l0bl1 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b1c341 l0bl1 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b1c342 l0bl1 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b1c343 l0bl1 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b1c344 l0bl1 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b1c345 l0bl1 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b1c346 l0bl1 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b1c347 l0bl1 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b1c348 l0bl1 vdd x348 x348b CELLD r1=10000e3 r0=900e3
xl0b1c349 l0bl1 vdd x349 x349b CELLD r1=10000e3 r0=900e3
xl0b1c350 l0bl1 vdd x350 x350b CELLD r1=10000e3 r0=900e3
xl0b1c351 l0bl1 vdd x351 x351b CELLD r1=10000e3 r0=900e3
xl0b1c352 l0bl1 vdd x352 x352b CELLD r1=10000e3 r0=900e3
xl0b1c353 l0bl1 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b1c354 l0bl1 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b1c355 l0bl1 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b1c356 l0bl1 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b1c357 l0bl1 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b1c358 l0bl1 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b1c359 l0bl1 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b1c360 l0bl1 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b1c361 l0bl1 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b1c362 l0bl1 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b1c363 l0bl1 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b1c364 l0bl1 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b1c365 l0bl1 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b1c366 l0bl1 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b1c367 l0bl1 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b1c368 l0bl1 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b1c369 l0bl1 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b1c370 l0bl1 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b1c371 l0bl1 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b1c372 l0bl1 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b1c373 l0bl1 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b1c374 l0bl1 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b1c375 l0bl1 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b1c376 l0bl1 vdd x376 x376b CELLD r1=10000e3 r0=900e3
xl0b1c377 l0bl1 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b1c378 l0bl1 vdd x378 x378b CELLD r1=10000e3 r0=900e3
xl0b1c379 l0bl1 vdd x379 x379b CELLD r1=10000e3 r0=900e3
xl0b1c380 l0bl1 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b1c381 l0bl1 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b1c382 l0bl1 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b1c383 l0bl1 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b1c384 l0bl1 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b1c385 l0bl1 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b1c386 l0bl1 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b1c387 l0bl1 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b1c388 l0bl1 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b1c389 l0bl1 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b1c390 l0bl1 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b1c391 l0bl1 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b1c392 l0bl1 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b1c393 l0bl1 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b1c394 l0bl1 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b1c395 l0bl1 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b1c396 l0bl1 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b1c397 l0bl1 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b1c398 l0bl1 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b1c399 l0bl1 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b1c400 l0bl1 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b1c401 l0bl1 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b1c402 l0bl1 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b1c403 l0bl1 vdd x403 x403b CELLD r1=10000e3 r0=900e3
xl0b1c404 l0bl1 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b1c405 l0bl1 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b1c406 l0bl1 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b1c407 l0bl1 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b1c408 l0bl1 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b1c409 l0bl1 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b1c410 l0bl1 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b1c411 l0bl1 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b1c412 l0bl1 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b1c413 l0bl1 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b1c414 l0bl1 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b1c415 l0bl1 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b1c416 l0bl1 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b1c417 l0bl1 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b1c418 l0bl1 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b1c419 l0bl1 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b1c420 l0bl1 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b1c421 l0bl1 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b1c422 l0bl1 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b1c423 l0bl1 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b1c424 l0bl1 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b1c425 l0bl1 vdd x425 x425b CELLD r1=900e3 r0=10000e3
xl0b1c426 l0bl1 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b1c427 l0bl1 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b1c428 l0bl1 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b1c429 l0bl1 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b1c430 l0bl1 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b1c431 l0bl1 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b1c432 l0bl1 vdd x432 x432b CELLD r1=10000e3 r0=900e3
xl0b1c433 l0bl1 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b1c434 l0bl1 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b1c435 l0bl1 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b1c436 l0bl1 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b1c437 l0bl1 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b1c438 l0bl1 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b1c439 l0bl1 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b1c440 l0bl1 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b1c441 l0bl1 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b1c442 l0bl1 vdd x442 x442b CELLD r1=900e3 r0=10000e3
xl0b1c443 l0bl1 vdd x443 x443b CELLD r1=900e3 r0=10000e3
xl0b1c444 l0bl1 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b1c445 l0bl1 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b1c446 l0bl1 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b1c447 l0bl1 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b1c448 l0bl1 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b1c449 l0bl1 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b1c450 l0bl1 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b1c451 l0bl1 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b1c452 l0bl1 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b1c453 l0bl1 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b1c454 l0bl1 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b1c455 l0bl1 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b1c456 l0bl1 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b1c457 l0bl1 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b1c458 l0bl1 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b1c459 l0bl1 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b1c460 l0bl1 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b1c461 l0bl1 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b1c462 l0bl1 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b1c463 l0bl1 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b1c464 l0bl1 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b1c465 l0bl1 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b1c466 l0bl1 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b1c467 l0bl1 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b1c468 l0bl1 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b1c469 l0bl1 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b1c470 l0bl1 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b1c471 l0bl1 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b1c472 l0bl1 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b1c473 l0bl1 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b1c474 l0bl1 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b1c475 l0bl1 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b1c476 l0bl1 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b1c477 l0bl1 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b1c478 l0bl1 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b1c479 l0bl1 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b1c480 l0bl1 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b1c481 l0bl1 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b1c482 l0bl1 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b1c483 l0bl1 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b1c484 l0bl1 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b1c485 l0bl1 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b1c486 l0bl1 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b1c487 l0bl1 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b1c488 l0bl1 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b1c489 l0bl1 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b1c490 l0bl1 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b1c491 l0bl1 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b1c492 l0bl1 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b1c493 l0bl1 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b1c494 l0bl1 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b1c495 l0bl1 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b1c496 l0bl1 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b1c497 l0bl1 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b1c498 l0bl1 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b1c499 l0bl1 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b1c500 l0bl1 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b1c501 l0bl1 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b1c502 l0bl1 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b1c503 l0bl1 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b1c504 l0bl1 vdd x504 x504b CELLD r1=10000e3 r0=900e3
xl0b1c505 l0bl1 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b1c506 l0bl1 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b1c507 l0bl1 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b1c508 l0bl1 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b1c509 l0bl1 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b1c510 l0bl1 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b1c511 l0bl1 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b1c512 l0bl1 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b1c513 l0bl1 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b1c514 l0bl1 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b1c515 l0bl1 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b1c516 l0bl1 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b1c517 l0bl1 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b1c518 l0bl1 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b1c519 l0bl1 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b1c520 l0bl1 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b1c521 l0bl1 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b1c522 l0bl1 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b1c523 l0bl1 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b1c524 l0bl1 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b1c525 l0bl1 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b1c526 l0bl1 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b1c527 l0bl1 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b1c528 l0bl1 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b1c529 l0bl1 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b1c530 l0bl1 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b1c531 l0bl1 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b1c532 l0bl1 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b1c533 l0bl1 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b1c534 l0bl1 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b1c535 l0bl1 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b1c536 l0bl1 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b1c537 l0bl1 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b1c538 l0bl1 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b1c539 l0bl1 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b1c540 l0bl1 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b1c541 l0bl1 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b1c542 l0bl1 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b1c543 l0bl1 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b1c544 l0bl1 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b1c545 l0bl1 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b1c546 l0bl1 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b1c547 l0bl1 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b1c548 l0bl1 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b1c549 l0bl1 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b1c550 l0bl1 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b1c551 l0bl1 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b1c552 l0bl1 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b1c553 l0bl1 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b1c554 l0bl1 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b1c555 l0bl1 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b1c556 l0bl1 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b1c557 l0bl1 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b1c558 l0bl1 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b1c559 l0bl1 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b1c560 l0bl1 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b1c561 l0bl1 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b1c562 l0bl1 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b1c563 l0bl1 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b1c564 l0bl1 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b1c565 l0bl1 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b1c566 l0bl1 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b1c567 l0bl1 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b1c568 l0bl1 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b1c569 l0bl1 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b1c570 l0bl1 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b1c571 l0bl1 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b1c572 l0bl1 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b1c573 l0bl1 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b1c574 l0bl1 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b1c575 l0bl1 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b1c576 l0bl1 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b1c577 l0bl1 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b1c578 l0bl1 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b1c579 l0bl1 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b1c580 l0bl1 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b1c581 l0bl1 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b1c582 l0bl1 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b1c583 l0bl1 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b1c584 l0bl1 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b1c585 l0bl1 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b1c586 l0bl1 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b1c587 l0bl1 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b1c588 l0bl1 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b1c589 l0bl1 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b1c590 l0bl1 vdd x590 x590b CELLD r1=10000e3 r0=900e3
xl0b1c591 l0bl1 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b1c592 l0bl1 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b1c593 l0bl1 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b1c594 l0bl1 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b1c595 l0bl1 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b1c596 l0bl1 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b1c597 l0bl1 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b1c598 l0bl1 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b1c599 l0bl1 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b1c600 l0bl1 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b1c601 l0bl1 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b1c602 l0bl1 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b1c603 l0bl1 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b1c604 l0bl1 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b1c605 l0bl1 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b1c606 l0bl1 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b1c607 l0bl1 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b1c608 l0bl1 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b1c609 l0bl1 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b1c610 l0bl1 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b1c611 l0bl1 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b1c612 l0bl1 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b1c613 l0bl1 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b1c614 l0bl1 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b1c615 l0bl1 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b1c616 l0bl1 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b1c617 l0bl1 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b1c618 l0bl1 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b1c619 l0bl1 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b1c620 l0bl1 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b1c621 l0bl1 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b1c622 l0bl1 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b1c623 l0bl1 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b1c624 l0bl1 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b1c625 l0bl1 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b1c626 l0bl1 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b1c627 l0bl1 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b1c628 l0bl1 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b1c629 l0bl1 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b1c630 l0bl1 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b1c631 l0bl1 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b1c632 l0bl1 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b1c633 l0bl1 vdd x633 x633b CELLD r1=10000e3 r0=900e3
xl0b1c634 l0bl1 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b1c635 l0bl1 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b1c636 l0bl1 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b1c637 l0bl1 vdd x637 x637b CELLD r1=10000e3 r0=900e3
xl0b1c638 l0bl1 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b1c639 l0bl1 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b1c640 l0bl1 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b1c641 l0bl1 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b1c642 l0bl1 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b1c643 l0bl1 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b1c644 l0bl1 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b1c645 l0bl1 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b1c646 l0bl1 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b1c647 l0bl1 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b1c648 l0bl1 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b1c649 l0bl1 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b1c650 l0bl1 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b1c651 l0bl1 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b1c652 l0bl1 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b1c653 l0bl1 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b1c654 l0bl1 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b1c655 l0bl1 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b1c656 l0bl1 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b1c657 l0bl1 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b1c658 l0bl1 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b1c659 l0bl1 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b1c660 l0bl1 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b1c661 l0bl1 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b1c662 l0bl1 vdd x662 x662b CELLD r1=10000e3 r0=900e3
xl0b1c663 l0bl1 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b1c664 l0bl1 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b1c665 l0bl1 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b1c666 l0bl1 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b1c667 l0bl1 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b1c668 l0bl1 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b1c669 l0bl1 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b1c670 l0bl1 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b1c671 l0bl1 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b1c672 l0bl1 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b1c673 l0bl1 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b1c674 l0bl1 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b1c675 l0bl1 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b1c676 l0bl1 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b1c677 l0bl1 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b1c678 l0bl1 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b1c679 l0bl1 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b1c680 l0bl1 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b1c681 l0bl1 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b1c682 l0bl1 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b1c683 l0bl1 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b1c684 l0bl1 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b1c685 l0bl1 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b1c686 l0bl1 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b1c687 l0bl1 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b1c688 l0bl1 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b1c689 l0bl1 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b1c690 l0bl1 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b1c691 l0bl1 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b1c692 l0bl1 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b1c693 l0bl1 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b1c694 l0bl1 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b1c695 l0bl1 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b1c696 l0bl1 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b1c697 l0bl1 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b1c698 l0bl1 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b1c699 l0bl1 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b1c700 l0bl1 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b1c701 l0bl1 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b1c702 l0bl1 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b1c703 l0bl1 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b1c704 l0bl1 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b1c705 l0bl1 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b1c706 l0bl1 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b1c707 l0bl1 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b1c708 l0bl1 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b1c709 l0bl1 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b1c710 l0bl1 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b1c711 l0bl1 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b1c712 l0bl1 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b1c713 l0bl1 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b1c714 l0bl1 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b1c715 l0bl1 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b1c716 l0bl1 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b1c717 l0bl1 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b1c718 l0bl1 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b1c719 l0bl1 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b1c720 l0bl1 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b1c721 l0bl1 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b1c722 l0bl1 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b1c723 l0bl1 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b1c724 l0bl1 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b1c725 l0bl1 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b1c726 l0bl1 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b1c727 l0bl1 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b1c728 l0bl1 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b1c729 l0bl1 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b1c730 l0bl1 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b1c731 l0bl1 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b1c732 l0bl1 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b1c733 l0bl1 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b1c734 l0bl1 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b1c735 l0bl1 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b1c736 l0bl1 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b1c737 l0bl1 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b1c738 l0bl1 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b1c739 l0bl1 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b1c740 l0bl1 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b1c741 l0bl1 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b1c742 l0bl1 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b1c743 l0bl1 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b1c744 l0bl1 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b1c745 l0bl1 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b1c746 l0bl1 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b1c747 l0bl1 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b1c748 l0bl1 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b1c749 l0bl1 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b1c750 l0bl1 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b1c751 l0bl1 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b1c752 l0bl1 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b1c753 l0bl1 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b1c754 l0bl1 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b1c755 l0bl1 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b1c756 l0bl1 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b1c757 l0bl1 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b1c758 l0bl1 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b1c759 l0bl1 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b1c760 l0bl1 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b1c761 l0bl1 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b1c762 l0bl1 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b1c763 l0bl1 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b1c764 l0bl1 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b1c765 l0bl1 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b1c766 l0bl1 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b1c767 l0bl1 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b1c768 l0bl1 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b1c769 l0bl1 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b1c770 l0bl1 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b1c771 l0bl1 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b1c772 l0bl1 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b1c773 l0bl1 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b1c774 l0bl1 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b1c775 l0bl1 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b1c776 l0bl1 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b1c777 l0bl1 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b1c778 l0bl1 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b1c779 l0bl1 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b1c780 l0bl1 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b1c781 l0bl1 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b1c782 l0bl1 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b1c783 l0bl1 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b2c0 l0bl2 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b2c1 l0bl2 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b2c2 l0bl2 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b2c3 l0bl2 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b2c4 l0bl2 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b2c5 l0bl2 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b2c6 l0bl2 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b2c7 l0bl2 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b2c8 l0bl2 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b2c9 l0bl2 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b2c10 l0bl2 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b2c11 l0bl2 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b2c12 l0bl2 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b2c13 l0bl2 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b2c14 l0bl2 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b2c15 l0bl2 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b2c16 l0bl2 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b2c17 l0bl2 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b2c18 l0bl2 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b2c19 l0bl2 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b2c20 l0bl2 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b2c21 l0bl2 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b2c22 l0bl2 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b2c23 l0bl2 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b2c24 l0bl2 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b2c25 l0bl2 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b2c26 l0bl2 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b2c27 l0bl2 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b2c28 l0bl2 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b2c29 l0bl2 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b2c30 l0bl2 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b2c31 l0bl2 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b2c32 l0bl2 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b2c33 l0bl2 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b2c34 l0bl2 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b2c35 l0bl2 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b2c36 l0bl2 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b2c37 l0bl2 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b2c38 l0bl2 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b2c39 l0bl2 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b2c40 l0bl2 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b2c41 l0bl2 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b2c42 l0bl2 vdd x42 x42b CELLD r1=10000e3 r0=900e3
xl0b2c43 l0bl2 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b2c44 l0bl2 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b2c45 l0bl2 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b2c46 l0bl2 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b2c47 l0bl2 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b2c48 l0bl2 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b2c49 l0bl2 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b2c50 l0bl2 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b2c51 l0bl2 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b2c52 l0bl2 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b2c53 l0bl2 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b2c54 l0bl2 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b2c55 l0bl2 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b2c56 l0bl2 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b2c57 l0bl2 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b2c58 l0bl2 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b2c59 l0bl2 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b2c60 l0bl2 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b2c61 l0bl2 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b2c62 l0bl2 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b2c63 l0bl2 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b2c64 l0bl2 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b2c65 l0bl2 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b2c66 l0bl2 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b2c67 l0bl2 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b2c68 l0bl2 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b2c69 l0bl2 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b2c70 l0bl2 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b2c71 l0bl2 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b2c72 l0bl2 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b2c73 l0bl2 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b2c74 l0bl2 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b2c75 l0bl2 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b2c76 l0bl2 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b2c77 l0bl2 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b2c78 l0bl2 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b2c79 l0bl2 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b2c80 l0bl2 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b2c81 l0bl2 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b2c82 l0bl2 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b2c83 l0bl2 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b2c84 l0bl2 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b2c85 l0bl2 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b2c86 l0bl2 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b2c87 l0bl2 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b2c88 l0bl2 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b2c89 l0bl2 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b2c90 l0bl2 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b2c91 l0bl2 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b2c92 l0bl2 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b2c93 l0bl2 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b2c94 l0bl2 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b2c95 l0bl2 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b2c96 l0bl2 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b2c97 l0bl2 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b2c98 l0bl2 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b2c99 l0bl2 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b2c100 l0bl2 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b2c101 l0bl2 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b2c102 l0bl2 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b2c103 l0bl2 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b2c104 l0bl2 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b2c105 l0bl2 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b2c106 l0bl2 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b2c107 l0bl2 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b2c108 l0bl2 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b2c109 l0bl2 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b2c110 l0bl2 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b2c111 l0bl2 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b2c112 l0bl2 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b2c113 l0bl2 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b2c114 l0bl2 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b2c115 l0bl2 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b2c116 l0bl2 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b2c117 l0bl2 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b2c118 l0bl2 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b2c119 l0bl2 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b2c120 l0bl2 vdd x120 x120b CELLD r1=900e3 r0=10000e3
xl0b2c121 l0bl2 vdd x121 x121b CELLD r1=900e3 r0=10000e3
xl0b2c122 l0bl2 vdd x122 x122b CELLD r1=900e3 r0=10000e3
xl0b2c123 l0bl2 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b2c124 l0bl2 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b2c125 l0bl2 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b2c126 l0bl2 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b2c127 l0bl2 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b2c128 l0bl2 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b2c129 l0bl2 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b2c130 l0bl2 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b2c131 l0bl2 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b2c132 l0bl2 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b2c133 l0bl2 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b2c134 l0bl2 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b2c135 l0bl2 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b2c136 l0bl2 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b2c137 l0bl2 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b2c138 l0bl2 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b2c139 l0bl2 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b2c140 l0bl2 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b2c141 l0bl2 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b2c142 l0bl2 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b2c143 l0bl2 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b2c144 l0bl2 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b2c145 l0bl2 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b2c146 l0bl2 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b2c147 l0bl2 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b2c148 l0bl2 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b2c149 l0bl2 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b2c150 l0bl2 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b2c151 l0bl2 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b2c152 l0bl2 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b2c153 l0bl2 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b2c154 l0bl2 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b2c155 l0bl2 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b2c156 l0bl2 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b2c157 l0bl2 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b2c158 l0bl2 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b2c159 l0bl2 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b2c160 l0bl2 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b2c161 l0bl2 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b2c162 l0bl2 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b2c163 l0bl2 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b2c164 l0bl2 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b2c165 l0bl2 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b2c166 l0bl2 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b2c167 l0bl2 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b2c168 l0bl2 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b2c169 l0bl2 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b2c170 l0bl2 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b2c171 l0bl2 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b2c172 l0bl2 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b2c173 l0bl2 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b2c174 l0bl2 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b2c175 l0bl2 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b2c176 l0bl2 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b2c177 l0bl2 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b2c178 l0bl2 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b2c179 l0bl2 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b2c180 l0bl2 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b2c181 l0bl2 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b2c182 l0bl2 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b2c183 l0bl2 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b2c184 l0bl2 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b2c185 l0bl2 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b2c186 l0bl2 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b2c187 l0bl2 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b2c188 l0bl2 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b2c189 l0bl2 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b2c190 l0bl2 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b2c191 l0bl2 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b2c192 l0bl2 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b2c193 l0bl2 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b2c194 l0bl2 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b2c195 l0bl2 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b2c196 l0bl2 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b2c197 l0bl2 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b2c198 l0bl2 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b2c199 l0bl2 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b2c200 l0bl2 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b2c201 l0bl2 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b2c202 l0bl2 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b2c203 l0bl2 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b2c204 l0bl2 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b2c205 l0bl2 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b2c206 l0bl2 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b2c207 l0bl2 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b2c208 l0bl2 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b2c209 l0bl2 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b2c210 l0bl2 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b2c211 l0bl2 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b2c212 l0bl2 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b2c213 l0bl2 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b2c214 l0bl2 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b2c215 l0bl2 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b2c216 l0bl2 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b2c217 l0bl2 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b2c218 l0bl2 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b2c219 l0bl2 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b2c220 l0bl2 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b2c221 l0bl2 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b2c222 l0bl2 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b2c223 l0bl2 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b2c224 l0bl2 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b2c225 l0bl2 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b2c226 l0bl2 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b2c227 l0bl2 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b2c228 l0bl2 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b2c229 l0bl2 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b2c230 l0bl2 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b2c231 l0bl2 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b2c232 l0bl2 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b2c233 l0bl2 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b2c234 l0bl2 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b2c235 l0bl2 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b2c236 l0bl2 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b2c237 l0bl2 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b2c238 l0bl2 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b2c239 l0bl2 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b2c240 l0bl2 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b2c241 l0bl2 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b2c242 l0bl2 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b2c243 l0bl2 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b2c244 l0bl2 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b2c245 l0bl2 vdd x245 x245b CELLD r1=900e3 r0=10000e3
xl0b2c246 l0bl2 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b2c247 l0bl2 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b2c248 l0bl2 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b2c249 l0bl2 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b2c250 l0bl2 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b2c251 l0bl2 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b2c252 l0bl2 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b2c253 l0bl2 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b2c254 l0bl2 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b2c255 l0bl2 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b2c256 l0bl2 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b2c257 l0bl2 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b2c258 l0bl2 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b2c259 l0bl2 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b2c260 l0bl2 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b2c261 l0bl2 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b2c262 l0bl2 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b2c263 l0bl2 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b2c264 l0bl2 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b2c265 l0bl2 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b2c266 l0bl2 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b2c267 l0bl2 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b2c268 l0bl2 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b2c269 l0bl2 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b2c270 l0bl2 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b2c271 l0bl2 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b2c272 l0bl2 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b2c273 l0bl2 vdd x273 x273b CELLD r1=900e3 r0=10000e3
xl0b2c274 l0bl2 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b2c275 l0bl2 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b2c276 l0bl2 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b2c277 l0bl2 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b2c278 l0bl2 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b2c279 l0bl2 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b2c280 l0bl2 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b2c281 l0bl2 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b2c282 l0bl2 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b2c283 l0bl2 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b2c284 l0bl2 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b2c285 l0bl2 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b2c286 l0bl2 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b2c287 l0bl2 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b2c288 l0bl2 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b2c289 l0bl2 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b2c290 l0bl2 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b2c291 l0bl2 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b2c292 l0bl2 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b2c293 l0bl2 vdd x293 x293b CELLD r1=900e3 r0=10000e3
xl0b2c294 l0bl2 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b2c295 l0bl2 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b2c296 l0bl2 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b2c297 l0bl2 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b2c298 l0bl2 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b2c299 l0bl2 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b2c300 l0bl2 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b2c301 l0bl2 vdd x301 x301b CELLD r1=900e3 r0=10000e3
xl0b2c302 l0bl2 vdd x302 x302b CELLD r1=900e3 r0=10000e3
xl0b2c303 l0bl2 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b2c304 l0bl2 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b2c305 l0bl2 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b2c306 l0bl2 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b2c307 l0bl2 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b2c308 l0bl2 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b2c309 l0bl2 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b2c310 l0bl2 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b2c311 l0bl2 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b2c312 l0bl2 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b2c313 l0bl2 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b2c314 l0bl2 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b2c315 l0bl2 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b2c316 l0bl2 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b2c317 l0bl2 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b2c318 l0bl2 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b2c319 l0bl2 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b2c320 l0bl2 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b2c321 l0bl2 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b2c322 l0bl2 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b2c323 l0bl2 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b2c324 l0bl2 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b2c325 l0bl2 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b2c326 l0bl2 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b2c327 l0bl2 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b2c328 l0bl2 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b2c329 l0bl2 vdd x329 x329b CELLD r1=900e3 r0=10000e3
xl0b2c330 l0bl2 vdd x330 x330b CELLD r1=900e3 r0=10000e3
xl0b2c331 l0bl2 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b2c332 l0bl2 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b2c333 l0bl2 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b2c334 l0bl2 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b2c335 l0bl2 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b2c336 l0bl2 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b2c337 l0bl2 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b2c338 l0bl2 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b2c339 l0bl2 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b2c340 l0bl2 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b2c341 l0bl2 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b2c342 l0bl2 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b2c343 l0bl2 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b2c344 l0bl2 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b2c345 l0bl2 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b2c346 l0bl2 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b2c347 l0bl2 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b2c348 l0bl2 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b2c349 l0bl2 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b2c350 l0bl2 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b2c351 l0bl2 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b2c352 l0bl2 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b2c353 l0bl2 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b2c354 l0bl2 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b2c355 l0bl2 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b2c356 l0bl2 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b2c357 l0bl2 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b2c358 l0bl2 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b2c359 l0bl2 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b2c360 l0bl2 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b2c361 l0bl2 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b2c362 l0bl2 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b2c363 l0bl2 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b2c364 l0bl2 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b2c365 l0bl2 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b2c366 l0bl2 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b2c367 l0bl2 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b2c368 l0bl2 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b2c369 l0bl2 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b2c370 l0bl2 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b2c371 l0bl2 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b2c372 l0bl2 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b2c373 l0bl2 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b2c374 l0bl2 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b2c375 l0bl2 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b2c376 l0bl2 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b2c377 l0bl2 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b2c378 l0bl2 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b2c379 l0bl2 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b2c380 l0bl2 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b2c381 l0bl2 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b2c382 l0bl2 vdd x382 x382b CELLD r1=10000e3 r0=900e3
xl0b2c383 l0bl2 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b2c384 l0bl2 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b2c385 l0bl2 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b2c386 l0bl2 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b2c387 l0bl2 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b2c388 l0bl2 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b2c389 l0bl2 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b2c390 l0bl2 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b2c391 l0bl2 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b2c392 l0bl2 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b2c393 l0bl2 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b2c394 l0bl2 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b2c395 l0bl2 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b2c396 l0bl2 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b2c397 l0bl2 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b2c398 l0bl2 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b2c399 l0bl2 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b2c400 l0bl2 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b2c401 l0bl2 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b2c402 l0bl2 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b2c403 l0bl2 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b2c404 l0bl2 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b2c405 l0bl2 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b2c406 l0bl2 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b2c407 l0bl2 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b2c408 l0bl2 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b2c409 l0bl2 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b2c410 l0bl2 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b2c411 l0bl2 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b2c412 l0bl2 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b2c413 l0bl2 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b2c414 l0bl2 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b2c415 l0bl2 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b2c416 l0bl2 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b2c417 l0bl2 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b2c418 l0bl2 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b2c419 l0bl2 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b2c420 l0bl2 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b2c421 l0bl2 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b2c422 l0bl2 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b2c423 l0bl2 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b2c424 l0bl2 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b2c425 l0bl2 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b2c426 l0bl2 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b2c427 l0bl2 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b2c428 l0bl2 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b2c429 l0bl2 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b2c430 l0bl2 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b2c431 l0bl2 vdd x431 x431b CELLD r1=10000e3 r0=900e3
xl0b2c432 l0bl2 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b2c433 l0bl2 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b2c434 l0bl2 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b2c435 l0bl2 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b2c436 l0bl2 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b2c437 l0bl2 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b2c438 l0bl2 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b2c439 l0bl2 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b2c440 l0bl2 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b2c441 l0bl2 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b2c442 l0bl2 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b2c443 l0bl2 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b2c444 l0bl2 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b2c445 l0bl2 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b2c446 l0bl2 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b2c447 l0bl2 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b2c448 l0bl2 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b2c449 l0bl2 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b2c450 l0bl2 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b2c451 l0bl2 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b2c452 l0bl2 vdd x452 x452b CELLD r1=900e3 r0=10000e3
xl0b2c453 l0bl2 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b2c454 l0bl2 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b2c455 l0bl2 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b2c456 l0bl2 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b2c457 l0bl2 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b2c458 l0bl2 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b2c459 l0bl2 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b2c460 l0bl2 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b2c461 l0bl2 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b2c462 l0bl2 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b2c463 l0bl2 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b2c464 l0bl2 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b2c465 l0bl2 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b2c466 l0bl2 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b2c467 l0bl2 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b2c468 l0bl2 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b2c469 l0bl2 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b2c470 l0bl2 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b2c471 l0bl2 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b2c472 l0bl2 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b2c473 l0bl2 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b2c474 l0bl2 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b2c475 l0bl2 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b2c476 l0bl2 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b2c477 l0bl2 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b2c478 l0bl2 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b2c479 l0bl2 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b2c480 l0bl2 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b2c481 l0bl2 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b2c482 l0bl2 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b2c483 l0bl2 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b2c484 l0bl2 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b2c485 l0bl2 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b2c486 l0bl2 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b2c487 l0bl2 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b2c488 l0bl2 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b2c489 l0bl2 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b2c490 l0bl2 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b2c491 l0bl2 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b2c492 l0bl2 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b2c493 l0bl2 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b2c494 l0bl2 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b2c495 l0bl2 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b2c496 l0bl2 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b2c497 l0bl2 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b2c498 l0bl2 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b2c499 l0bl2 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b2c500 l0bl2 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b2c501 l0bl2 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b2c502 l0bl2 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b2c503 l0bl2 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b2c504 l0bl2 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b2c505 l0bl2 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b2c506 l0bl2 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b2c507 l0bl2 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b2c508 l0bl2 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b2c509 l0bl2 vdd x509 x509b CELLD r1=900e3 r0=10000e3
xl0b2c510 l0bl2 vdd x510 x510b CELLD r1=900e3 r0=10000e3
xl0b2c511 l0bl2 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b2c512 l0bl2 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b2c513 l0bl2 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b2c514 l0bl2 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b2c515 l0bl2 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b2c516 l0bl2 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b2c517 l0bl2 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b2c518 l0bl2 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b2c519 l0bl2 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b2c520 l0bl2 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b2c521 l0bl2 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b2c522 l0bl2 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b2c523 l0bl2 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b2c524 l0bl2 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b2c525 l0bl2 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b2c526 l0bl2 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b2c527 l0bl2 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b2c528 l0bl2 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b2c529 l0bl2 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b2c530 l0bl2 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b2c531 l0bl2 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b2c532 l0bl2 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b2c533 l0bl2 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b2c534 l0bl2 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b2c535 l0bl2 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b2c536 l0bl2 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b2c537 l0bl2 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b2c538 l0bl2 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b2c539 l0bl2 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b2c540 l0bl2 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b2c541 l0bl2 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b2c542 l0bl2 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b2c543 l0bl2 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b2c544 l0bl2 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b2c545 l0bl2 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b2c546 l0bl2 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b2c547 l0bl2 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b2c548 l0bl2 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b2c549 l0bl2 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b2c550 l0bl2 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b2c551 l0bl2 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b2c552 l0bl2 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b2c553 l0bl2 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b2c554 l0bl2 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b2c555 l0bl2 vdd x555 x555b CELLD r1=900e3 r0=10000e3
xl0b2c556 l0bl2 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b2c557 l0bl2 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b2c558 l0bl2 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b2c559 l0bl2 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b2c560 l0bl2 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b2c561 l0bl2 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b2c562 l0bl2 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b2c563 l0bl2 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b2c564 l0bl2 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b2c565 l0bl2 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b2c566 l0bl2 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b2c567 l0bl2 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b2c568 l0bl2 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b2c569 l0bl2 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b2c570 l0bl2 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b2c571 l0bl2 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b2c572 l0bl2 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b2c573 l0bl2 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b2c574 l0bl2 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b2c575 l0bl2 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b2c576 l0bl2 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b2c577 l0bl2 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b2c578 l0bl2 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b2c579 l0bl2 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b2c580 l0bl2 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b2c581 l0bl2 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b2c582 l0bl2 vdd x582 x582b CELLD r1=900e3 r0=10000e3
xl0b2c583 l0bl2 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b2c584 l0bl2 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b2c585 l0bl2 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b2c586 l0bl2 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b2c587 l0bl2 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b2c588 l0bl2 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b2c589 l0bl2 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b2c590 l0bl2 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b2c591 l0bl2 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b2c592 l0bl2 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b2c593 l0bl2 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b2c594 l0bl2 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b2c595 l0bl2 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b2c596 l0bl2 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b2c597 l0bl2 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b2c598 l0bl2 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b2c599 l0bl2 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b2c600 l0bl2 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b2c601 l0bl2 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b2c602 l0bl2 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b2c603 l0bl2 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b2c604 l0bl2 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b2c605 l0bl2 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b2c606 l0bl2 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b2c607 l0bl2 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b2c608 l0bl2 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b2c609 l0bl2 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b2c610 l0bl2 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b2c611 l0bl2 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b2c612 l0bl2 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b2c613 l0bl2 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b2c614 l0bl2 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b2c615 l0bl2 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b2c616 l0bl2 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b2c617 l0bl2 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b2c618 l0bl2 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b2c619 l0bl2 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b2c620 l0bl2 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b2c621 l0bl2 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b2c622 l0bl2 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b2c623 l0bl2 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b2c624 l0bl2 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b2c625 l0bl2 vdd x625 x625b CELLD r1=900e3 r0=10000e3
xl0b2c626 l0bl2 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b2c627 l0bl2 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b2c628 l0bl2 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b2c629 l0bl2 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b2c630 l0bl2 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b2c631 l0bl2 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b2c632 l0bl2 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b2c633 l0bl2 vdd x633 x633b CELLD r1=10000e3 r0=900e3
xl0b2c634 l0bl2 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b2c635 l0bl2 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b2c636 l0bl2 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b2c637 l0bl2 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b2c638 l0bl2 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b2c639 l0bl2 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b2c640 l0bl2 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b2c641 l0bl2 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b2c642 l0bl2 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b2c643 l0bl2 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b2c644 l0bl2 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b2c645 l0bl2 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b2c646 l0bl2 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b2c647 l0bl2 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b2c648 l0bl2 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b2c649 l0bl2 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b2c650 l0bl2 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b2c651 l0bl2 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b2c652 l0bl2 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b2c653 l0bl2 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b2c654 l0bl2 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b2c655 l0bl2 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b2c656 l0bl2 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b2c657 l0bl2 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b2c658 l0bl2 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b2c659 l0bl2 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b2c660 l0bl2 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b2c661 l0bl2 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b2c662 l0bl2 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b2c663 l0bl2 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b2c664 l0bl2 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b2c665 l0bl2 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b2c666 l0bl2 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b2c667 l0bl2 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b2c668 l0bl2 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b2c669 l0bl2 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b2c670 l0bl2 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b2c671 l0bl2 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b2c672 l0bl2 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b2c673 l0bl2 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b2c674 l0bl2 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b2c675 l0bl2 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b2c676 l0bl2 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b2c677 l0bl2 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b2c678 l0bl2 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b2c679 l0bl2 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b2c680 l0bl2 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b2c681 l0bl2 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b2c682 l0bl2 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b2c683 l0bl2 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b2c684 l0bl2 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b2c685 l0bl2 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b2c686 l0bl2 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b2c687 l0bl2 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b2c688 l0bl2 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b2c689 l0bl2 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b2c690 l0bl2 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b2c691 l0bl2 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b2c692 l0bl2 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b2c693 l0bl2 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b2c694 l0bl2 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b2c695 l0bl2 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b2c696 l0bl2 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b2c697 l0bl2 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b2c698 l0bl2 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b2c699 l0bl2 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b2c700 l0bl2 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b2c701 l0bl2 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b2c702 l0bl2 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b2c703 l0bl2 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b2c704 l0bl2 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b2c705 l0bl2 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b2c706 l0bl2 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b2c707 l0bl2 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b2c708 l0bl2 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b2c709 l0bl2 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b2c710 l0bl2 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b2c711 l0bl2 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b2c712 l0bl2 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b2c713 l0bl2 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b2c714 l0bl2 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b2c715 l0bl2 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b2c716 l0bl2 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b2c717 l0bl2 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b2c718 l0bl2 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b2c719 l0bl2 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b2c720 l0bl2 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b2c721 l0bl2 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b2c722 l0bl2 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b2c723 l0bl2 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b2c724 l0bl2 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b2c725 l0bl2 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b2c726 l0bl2 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b2c727 l0bl2 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b2c728 l0bl2 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b2c729 l0bl2 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b2c730 l0bl2 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b2c731 l0bl2 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b2c732 l0bl2 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b2c733 l0bl2 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b2c734 l0bl2 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b2c735 l0bl2 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b2c736 l0bl2 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b2c737 l0bl2 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b2c738 l0bl2 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b2c739 l0bl2 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b2c740 l0bl2 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b2c741 l0bl2 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b2c742 l0bl2 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b2c743 l0bl2 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b2c744 l0bl2 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b2c745 l0bl2 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b2c746 l0bl2 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b2c747 l0bl2 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b2c748 l0bl2 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b2c749 l0bl2 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b2c750 l0bl2 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b2c751 l0bl2 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b2c752 l0bl2 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b2c753 l0bl2 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b2c754 l0bl2 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b2c755 l0bl2 vdd x755 x755b CELLD r1=10000e3 r0=900e3
xl0b2c756 l0bl2 vdd x756 x756b CELLD r1=900e3 r0=10000e3
xl0b2c757 l0bl2 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b2c758 l0bl2 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b2c759 l0bl2 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b2c760 l0bl2 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b2c761 l0bl2 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b2c762 l0bl2 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b2c763 l0bl2 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b2c764 l0bl2 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b2c765 l0bl2 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b2c766 l0bl2 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b2c767 l0bl2 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b2c768 l0bl2 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b2c769 l0bl2 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b2c770 l0bl2 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b2c771 l0bl2 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b2c772 l0bl2 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b2c773 l0bl2 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b2c774 l0bl2 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b2c775 l0bl2 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b2c776 l0bl2 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b2c777 l0bl2 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b2c778 l0bl2 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b2c779 l0bl2 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b2c780 l0bl2 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b2c781 l0bl2 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b2c782 l0bl2 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b2c783 l0bl2 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b3c0 l0bl3 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b3c1 l0bl3 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b3c2 l0bl3 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b3c3 l0bl3 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b3c4 l0bl3 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b3c5 l0bl3 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b3c6 l0bl3 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b3c7 l0bl3 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b3c8 l0bl3 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b3c9 l0bl3 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b3c10 l0bl3 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b3c11 l0bl3 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b3c12 l0bl3 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b3c13 l0bl3 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b3c14 l0bl3 vdd x14 x14b CELLD r1=10000e3 r0=900e3
xl0b3c15 l0bl3 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b3c16 l0bl3 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b3c17 l0bl3 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b3c18 l0bl3 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b3c19 l0bl3 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b3c20 l0bl3 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b3c21 l0bl3 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b3c22 l0bl3 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b3c23 l0bl3 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b3c24 l0bl3 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b3c25 l0bl3 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b3c26 l0bl3 vdd x26 x26b CELLD r1=10000e3 r0=900e3
xl0b3c27 l0bl3 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b3c28 l0bl3 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b3c29 l0bl3 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b3c30 l0bl3 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b3c31 l0bl3 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b3c32 l0bl3 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b3c33 l0bl3 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b3c34 l0bl3 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b3c35 l0bl3 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b3c36 l0bl3 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b3c37 l0bl3 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b3c38 l0bl3 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b3c39 l0bl3 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b3c40 l0bl3 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b3c41 l0bl3 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b3c42 l0bl3 vdd x42 x42b CELLD r1=10000e3 r0=900e3
xl0b3c43 l0bl3 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b3c44 l0bl3 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b3c45 l0bl3 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b3c46 l0bl3 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b3c47 l0bl3 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b3c48 l0bl3 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b3c49 l0bl3 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b3c50 l0bl3 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b3c51 l0bl3 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b3c52 l0bl3 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b3c53 l0bl3 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b3c54 l0bl3 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b3c55 l0bl3 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b3c56 l0bl3 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b3c57 l0bl3 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b3c58 l0bl3 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b3c59 l0bl3 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b3c60 l0bl3 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b3c61 l0bl3 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b3c62 l0bl3 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b3c63 l0bl3 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b3c64 l0bl3 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b3c65 l0bl3 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b3c66 l0bl3 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b3c67 l0bl3 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b3c68 l0bl3 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b3c69 l0bl3 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b3c70 l0bl3 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b3c71 l0bl3 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b3c72 l0bl3 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b3c73 l0bl3 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b3c74 l0bl3 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b3c75 l0bl3 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b3c76 l0bl3 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b3c77 l0bl3 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b3c78 l0bl3 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b3c79 l0bl3 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b3c80 l0bl3 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b3c81 l0bl3 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b3c82 l0bl3 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b3c83 l0bl3 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b3c84 l0bl3 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b3c85 l0bl3 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b3c86 l0bl3 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b3c87 l0bl3 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b3c88 l0bl3 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b3c89 l0bl3 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b3c90 l0bl3 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b3c91 l0bl3 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b3c92 l0bl3 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b3c93 l0bl3 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b3c94 l0bl3 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b3c95 l0bl3 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b3c96 l0bl3 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b3c97 l0bl3 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b3c98 l0bl3 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b3c99 l0bl3 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b3c100 l0bl3 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b3c101 l0bl3 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b3c102 l0bl3 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b3c103 l0bl3 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b3c104 l0bl3 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b3c105 l0bl3 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b3c106 l0bl3 vdd x106 x106b CELLD r1=10000e3 r0=900e3
xl0b3c107 l0bl3 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b3c108 l0bl3 vdd x108 x108b CELLD r1=10000e3 r0=900e3
xl0b3c109 l0bl3 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b3c110 l0bl3 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b3c111 l0bl3 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b3c112 l0bl3 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b3c113 l0bl3 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b3c114 l0bl3 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b3c115 l0bl3 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b3c116 l0bl3 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b3c117 l0bl3 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b3c118 l0bl3 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b3c119 l0bl3 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b3c120 l0bl3 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b3c121 l0bl3 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b3c122 l0bl3 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b3c123 l0bl3 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b3c124 l0bl3 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b3c125 l0bl3 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b3c126 l0bl3 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b3c127 l0bl3 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b3c128 l0bl3 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b3c129 l0bl3 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b3c130 l0bl3 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b3c131 l0bl3 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b3c132 l0bl3 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b3c133 l0bl3 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b3c134 l0bl3 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b3c135 l0bl3 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b3c136 l0bl3 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b3c137 l0bl3 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b3c138 l0bl3 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b3c139 l0bl3 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b3c140 l0bl3 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b3c141 l0bl3 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b3c142 l0bl3 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b3c143 l0bl3 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b3c144 l0bl3 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b3c145 l0bl3 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b3c146 l0bl3 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b3c147 l0bl3 vdd x147 x147b CELLD r1=900e3 r0=10000e3
xl0b3c148 l0bl3 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b3c149 l0bl3 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b3c150 l0bl3 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b3c151 l0bl3 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b3c152 l0bl3 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b3c153 l0bl3 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b3c154 l0bl3 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b3c155 l0bl3 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b3c156 l0bl3 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b3c157 l0bl3 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b3c158 l0bl3 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b3c159 l0bl3 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b3c160 l0bl3 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b3c161 l0bl3 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b3c162 l0bl3 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b3c163 l0bl3 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b3c164 l0bl3 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b3c165 l0bl3 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b3c166 l0bl3 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b3c167 l0bl3 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b3c168 l0bl3 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b3c169 l0bl3 vdd x169 x169b CELLD r1=10000e3 r0=900e3
xl0b3c170 l0bl3 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b3c171 l0bl3 vdd x171 x171b CELLD r1=10000e3 r0=900e3
xl0b3c172 l0bl3 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b3c173 l0bl3 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b3c174 l0bl3 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b3c175 l0bl3 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b3c176 l0bl3 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b3c177 l0bl3 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b3c178 l0bl3 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b3c179 l0bl3 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b3c180 l0bl3 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b3c181 l0bl3 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b3c182 l0bl3 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b3c183 l0bl3 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b3c184 l0bl3 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b3c185 l0bl3 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b3c186 l0bl3 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b3c187 l0bl3 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b3c188 l0bl3 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b3c189 l0bl3 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b3c190 l0bl3 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b3c191 l0bl3 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b3c192 l0bl3 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b3c193 l0bl3 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b3c194 l0bl3 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b3c195 l0bl3 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b3c196 l0bl3 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b3c197 l0bl3 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b3c198 l0bl3 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b3c199 l0bl3 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b3c200 l0bl3 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b3c201 l0bl3 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b3c202 l0bl3 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b3c203 l0bl3 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b3c204 l0bl3 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b3c205 l0bl3 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b3c206 l0bl3 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b3c207 l0bl3 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b3c208 l0bl3 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b3c209 l0bl3 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b3c210 l0bl3 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b3c211 l0bl3 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b3c212 l0bl3 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b3c213 l0bl3 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b3c214 l0bl3 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b3c215 l0bl3 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b3c216 l0bl3 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b3c217 l0bl3 vdd x217 x217b CELLD r1=900e3 r0=10000e3
xl0b3c218 l0bl3 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b3c219 l0bl3 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b3c220 l0bl3 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b3c221 l0bl3 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b3c222 l0bl3 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b3c223 l0bl3 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b3c224 l0bl3 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b3c225 l0bl3 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b3c226 l0bl3 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b3c227 l0bl3 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b3c228 l0bl3 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b3c229 l0bl3 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b3c230 l0bl3 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b3c231 l0bl3 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b3c232 l0bl3 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b3c233 l0bl3 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b3c234 l0bl3 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b3c235 l0bl3 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b3c236 l0bl3 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b3c237 l0bl3 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b3c238 l0bl3 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b3c239 l0bl3 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b3c240 l0bl3 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b3c241 l0bl3 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b3c242 l0bl3 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b3c243 l0bl3 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b3c244 l0bl3 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b3c245 l0bl3 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b3c246 l0bl3 vdd x246 x246b CELLD r1=900e3 r0=10000e3
xl0b3c247 l0bl3 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b3c248 l0bl3 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b3c249 l0bl3 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b3c250 l0bl3 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b3c251 l0bl3 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b3c252 l0bl3 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b3c253 l0bl3 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b3c254 l0bl3 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b3c255 l0bl3 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b3c256 l0bl3 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b3c257 l0bl3 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b3c258 l0bl3 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b3c259 l0bl3 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b3c260 l0bl3 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b3c261 l0bl3 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b3c262 l0bl3 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b3c263 l0bl3 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b3c264 l0bl3 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b3c265 l0bl3 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b3c266 l0bl3 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b3c267 l0bl3 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b3c268 l0bl3 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b3c269 l0bl3 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b3c270 l0bl3 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b3c271 l0bl3 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b3c272 l0bl3 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b3c273 l0bl3 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b3c274 l0bl3 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b3c275 l0bl3 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b3c276 l0bl3 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b3c277 l0bl3 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b3c278 l0bl3 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b3c279 l0bl3 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b3c280 l0bl3 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b3c281 l0bl3 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b3c282 l0bl3 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b3c283 l0bl3 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b3c284 l0bl3 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b3c285 l0bl3 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b3c286 l0bl3 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b3c287 l0bl3 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b3c288 l0bl3 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b3c289 l0bl3 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b3c290 l0bl3 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b3c291 l0bl3 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b3c292 l0bl3 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b3c293 l0bl3 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b3c294 l0bl3 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b3c295 l0bl3 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b3c296 l0bl3 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b3c297 l0bl3 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b3c298 l0bl3 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b3c299 l0bl3 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b3c300 l0bl3 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b3c301 l0bl3 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b3c302 l0bl3 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b3c303 l0bl3 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b3c304 l0bl3 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b3c305 l0bl3 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b3c306 l0bl3 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b3c307 l0bl3 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b3c308 l0bl3 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b3c309 l0bl3 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b3c310 l0bl3 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b3c311 l0bl3 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b3c312 l0bl3 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b3c313 l0bl3 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b3c314 l0bl3 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b3c315 l0bl3 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b3c316 l0bl3 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b3c317 l0bl3 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b3c318 l0bl3 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b3c319 l0bl3 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b3c320 l0bl3 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b3c321 l0bl3 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b3c322 l0bl3 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b3c323 l0bl3 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b3c324 l0bl3 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b3c325 l0bl3 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b3c326 l0bl3 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b3c327 l0bl3 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b3c328 l0bl3 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b3c329 l0bl3 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b3c330 l0bl3 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b3c331 l0bl3 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b3c332 l0bl3 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b3c333 l0bl3 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b3c334 l0bl3 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b3c335 l0bl3 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b3c336 l0bl3 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b3c337 l0bl3 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b3c338 l0bl3 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b3c339 l0bl3 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b3c340 l0bl3 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b3c341 l0bl3 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b3c342 l0bl3 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b3c343 l0bl3 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b3c344 l0bl3 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b3c345 l0bl3 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b3c346 l0bl3 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b3c347 l0bl3 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b3c348 l0bl3 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b3c349 l0bl3 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b3c350 l0bl3 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b3c351 l0bl3 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b3c352 l0bl3 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b3c353 l0bl3 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b3c354 l0bl3 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b3c355 l0bl3 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b3c356 l0bl3 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b3c357 l0bl3 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b3c358 l0bl3 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b3c359 l0bl3 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b3c360 l0bl3 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b3c361 l0bl3 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b3c362 l0bl3 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b3c363 l0bl3 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b3c364 l0bl3 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b3c365 l0bl3 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b3c366 l0bl3 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b3c367 l0bl3 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b3c368 l0bl3 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b3c369 l0bl3 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b3c370 l0bl3 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b3c371 l0bl3 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b3c372 l0bl3 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b3c373 l0bl3 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b3c374 l0bl3 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b3c375 l0bl3 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b3c376 l0bl3 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b3c377 l0bl3 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b3c378 l0bl3 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b3c379 l0bl3 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b3c380 l0bl3 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b3c381 l0bl3 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b3c382 l0bl3 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b3c383 l0bl3 vdd x383 x383b CELLD r1=10000e3 r0=900e3
xl0b3c384 l0bl3 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b3c385 l0bl3 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b3c386 l0bl3 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b3c387 l0bl3 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b3c388 l0bl3 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b3c389 l0bl3 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b3c390 l0bl3 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b3c391 l0bl3 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b3c392 l0bl3 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b3c393 l0bl3 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b3c394 l0bl3 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b3c395 l0bl3 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b3c396 l0bl3 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b3c397 l0bl3 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b3c398 l0bl3 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b3c399 l0bl3 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b3c400 l0bl3 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b3c401 l0bl3 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b3c402 l0bl3 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b3c403 l0bl3 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b3c404 l0bl3 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b3c405 l0bl3 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b3c406 l0bl3 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b3c407 l0bl3 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b3c408 l0bl3 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b3c409 l0bl3 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b3c410 l0bl3 vdd x410 x410b CELLD r1=10000e3 r0=900e3
xl0b3c411 l0bl3 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b3c412 l0bl3 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b3c413 l0bl3 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b3c414 l0bl3 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b3c415 l0bl3 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b3c416 l0bl3 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b3c417 l0bl3 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b3c418 l0bl3 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b3c419 l0bl3 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b3c420 l0bl3 vdd x420 x420b CELLD r1=10000e3 r0=900e3
xl0b3c421 l0bl3 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b3c422 l0bl3 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b3c423 l0bl3 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b3c424 l0bl3 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b3c425 l0bl3 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b3c426 l0bl3 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b3c427 l0bl3 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b3c428 l0bl3 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b3c429 l0bl3 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b3c430 l0bl3 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b3c431 l0bl3 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b3c432 l0bl3 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b3c433 l0bl3 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b3c434 l0bl3 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b3c435 l0bl3 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b3c436 l0bl3 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b3c437 l0bl3 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b3c438 l0bl3 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b3c439 l0bl3 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b3c440 l0bl3 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b3c441 l0bl3 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b3c442 l0bl3 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b3c443 l0bl3 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b3c444 l0bl3 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b3c445 l0bl3 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b3c446 l0bl3 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b3c447 l0bl3 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b3c448 l0bl3 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b3c449 l0bl3 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b3c450 l0bl3 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b3c451 l0bl3 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b3c452 l0bl3 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b3c453 l0bl3 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b3c454 l0bl3 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b3c455 l0bl3 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b3c456 l0bl3 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b3c457 l0bl3 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b3c458 l0bl3 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b3c459 l0bl3 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b3c460 l0bl3 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b3c461 l0bl3 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b3c462 l0bl3 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b3c463 l0bl3 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b3c464 l0bl3 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b3c465 l0bl3 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b3c466 l0bl3 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b3c467 l0bl3 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b3c468 l0bl3 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b3c469 l0bl3 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b3c470 l0bl3 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b3c471 l0bl3 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b3c472 l0bl3 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b3c473 l0bl3 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b3c474 l0bl3 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b3c475 l0bl3 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b3c476 l0bl3 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b3c477 l0bl3 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b3c478 l0bl3 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b3c479 l0bl3 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b3c480 l0bl3 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b3c481 l0bl3 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b3c482 l0bl3 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b3c483 l0bl3 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b3c484 l0bl3 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b3c485 l0bl3 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b3c486 l0bl3 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b3c487 l0bl3 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b3c488 l0bl3 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b3c489 l0bl3 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b3c490 l0bl3 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b3c491 l0bl3 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b3c492 l0bl3 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b3c493 l0bl3 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b3c494 l0bl3 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b3c495 l0bl3 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b3c496 l0bl3 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b3c497 l0bl3 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b3c498 l0bl3 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b3c499 l0bl3 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b3c500 l0bl3 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b3c501 l0bl3 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b3c502 l0bl3 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b3c503 l0bl3 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b3c504 l0bl3 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b3c505 l0bl3 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b3c506 l0bl3 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b3c507 l0bl3 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b3c508 l0bl3 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b3c509 l0bl3 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b3c510 l0bl3 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b3c511 l0bl3 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b3c512 l0bl3 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b3c513 l0bl3 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b3c514 l0bl3 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b3c515 l0bl3 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b3c516 l0bl3 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b3c517 l0bl3 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b3c518 l0bl3 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b3c519 l0bl3 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b3c520 l0bl3 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b3c521 l0bl3 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b3c522 l0bl3 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b3c523 l0bl3 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b3c524 l0bl3 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b3c525 l0bl3 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b3c526 l0bl3 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b3c527 l0bl3 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b3c528 l0bl3 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b3c529 l0bl3 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b3c530 l0bl3 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b3c531 l0bl3 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b3c532 l0bl3 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b3c533 l0bl3 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b3c534 l0bl3 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b3c535 l0bl3 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b3c536 l0bl3 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b3c537 l0bl3 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b3c538 l0bl3 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b3c539 l0bl3 vdd x539 x539b CELLD r1=900e3 r0=10000e3
xl0b3c540 l0bl3 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b3c541 l0bl3 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b3c542 l0bl3 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b3c543 l0bl3 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b3c544 l0bl3 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b3c545 l0bl3 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b3c546 l0bl3 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b3c547 l0bl3 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b3c548 l0bl3 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b3c549 l0bl3 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b3c550 l0bl3 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b3c551 l0bl3 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b3c552 l0bl3 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b3c553 l0bl3 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b3c554 l0bl3 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b3c555 l0bl3 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b3c556 l0bl3 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b3c557 l0bl3 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b3c558 l0bl3 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b3c559 l0bl3 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b3c560 l0bl3 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b3c561 l0bl3 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b3c562 l0bl3 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b3c563 l0bl3 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b3c564 l0bl3 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b3c565 l0bl3 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b3c566 l0bl3 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b3c567 l0bl3 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b3c568 l0bl3 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b3c569 l0bl3 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b3c570 l0bl3 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b3c571 l0bl3 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b3c572 l0bl3 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b3c573 l0bl3 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b3c574 l0bl3 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b3c575 l0bl3 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b3c576 l0bl3 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b3c577 l0bl3 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b3c578 l0bl3 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b3c579 l0bl3 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b3c580 l0bl3 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b3c581 l0bl3 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b3c582 l0bl3 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b3c583 l0bl3 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b3c584 l0bl3 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b3c585 l0bl3 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b3c586 l0bl3 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b3c587 l0bl3 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b3c588 l0bl3 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b3c589 l0bl3 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b3c590 l0bl3 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b3c591 l0bl3 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b3c592 l0bl3 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b3c593 l0bl3 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b3c594 l0bl3 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b3c595 l0bl3 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b3c596 l0bl3 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b3c597 l0bl3 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b3c598 l0bl3 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b3c599 l0bl3 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b3c600 l0bl3 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b3c601 l0bl3 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b3c602 l0bl3 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b3c603 l0bl3 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b3c604 l0bl3 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b3c605 l0bl3 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b3c606 l0bl3 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b3c607 l0bl3 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b3c608 l0bl3 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b3c609 l0bl3 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b3c610 l0bl3 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b3c611 l0bl3 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b3c612 l0bl3 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b3c613 l0bl3 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b3c614 l0bl3 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b3c615 l0bl3 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b3c616 l0bl3 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b3c617 l0bl3 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b3c618 l0bl3 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b3c619 l0bl3 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b3c620 l0bl3 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b3c621 l0bl3 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b3c622 l0bl3 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b3c623 l0bl3 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b3c624 l0bl3 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b3c625 l0bl3 vdd x625 x625b CELLD r1=900e3 r0=10000e3
xl0b3c626 l0bl3 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b3c627 l0bl3 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b3c628 l0bl3 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b3c629 l0bl3 vdd x629 x629b CELLD r1=900e3 r0=10000e3
xl0b3c630 l0bl3 vdd x630 x630b CELLD r1=900e3 r0=10000e3
xl0b3c631 l0bl3 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b3c632 l0bl3 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b3c633 l0bl3 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b3c634 l0bl3 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b3c635 l0bl3 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b3c636 l0bl3 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b3c637 l0bl3 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b3c638 l0bl3 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b3c639 l0bl3 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b3c640 l0bl3 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b3c641 l0bl3 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b3c642 l0bl3 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b3c643 l0bl3 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b3c644 l0bl3 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b3c645 l0bl3 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b3c646 l0bl3 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b3c647 l0bl3 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b3c648 l0bl3 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b3c649 l0bl3 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b3c650 l0bl3 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b3c651 l0bl3 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b3c652 l0bl3 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b3c653 l0bl3 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b3c654 l0bl3 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b3c655 l0bl3 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b3c656 l0bl3 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b3c657 l0bl3 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b3c658 l0bl3 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b3c659 l0bl3 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b3c660 l0bl3 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b3c661 l0bl3 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b3c662 l0bl3 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b3c663 l0bl3 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b3c664 l0bl3 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b3c665 l0bl3 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b3c666 l0bl3 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b3c667 l0bl3 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b3c668 l0bl3 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b3c669 l0bl3 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b3c670 l0bl3 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b3c671 l0bl3 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b3c672 l0bl3 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b3c673 l0bl3 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b3c674 l0bl3 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b3c675 l0bl3 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b3c676 l0bl3 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b3c677 l0bl3 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b3c678 l0bl3 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b3c679 l0bl3 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b3c680 l0bl3 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b3c681 l0bl3 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b3c682 l0bl3 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b3c683 l0bl3 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b3c684 l0bl3 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b3c685 l0bl3 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b3c686 l0bl3 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b3c687 l0bl3 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b3c688 l0bl3 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b3c689 l0bl3 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b3c690 l0bl3 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b3c691 l0bl3 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b3c692 l0bl3 vdd x692 x692b CELLD r1=10000e3 r0=900e3
xl0b3c693 l0bl3 vdd x693 x693b CELLD r1=10000e3 r0=900e3
xl0b3c694 l0bl3 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b3c695 l0bl3 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b3c696 l0bl3 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b3c697 l0bl3 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b3c698 l0bl3 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b3c699 l0bl3 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b3c700 l0bl3 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b3c701 l0bl3 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b3c702 l0bl3 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b3c703 l0bl3 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b3c704 l0bl3 vdd x704 x704b CELLD r1=10000e3 r0=900e3
xl0b3c705 l0bl3 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b3c706 l0bl3 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b3c707 l0bl3 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b3c708 l0bl3 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b3c709 l0bl3 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b3c710 l0bl3 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b3c711 l0bl3 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b3c712 l0bl3 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b3c713 l0bl3 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b3c714 l0bl3 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b3c715 l0bl3 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b3c716 l0bl3 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b3c717 l0bl3 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b3c718 l0bl3 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b3c719 l0bl3 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b3c720 l0bl3 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b3c721 l0bl3 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b3c722 l0bl3 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b3c723 l0bl3 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b3c724 l0bl3 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b3c725 l0bl3 vdd x725 x725b CELLD r1=10000e3 r0=900e3
xl0b3c726 l0bl3 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b3c727 l0bl3 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b3c728 l0bl3 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b3c729 l0bl3 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b3c730 l0bl3 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b3c731 l0bl3 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b3c732 l0bl3 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b3c733 l0bl3 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b3c734 l0bl3 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b3c735 l0bl3 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b3c736 l0bl3 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b3c737 l0bl3 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b3c738 l0bl3 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b3c739 l0bl3 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b3c740 l0bl3 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b3c741 l0bl3 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b3c742 l0bl3 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b3c743 l0bl3 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b3c744 l0bl3 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b3c745 l0bl3 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b3c746 l0bl3 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b3c747 l0bl3 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b3c748 l0bl3 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b3c749 l0bl3 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b3c750 l0bl3 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b3c751 l0bl3 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b3c752 l0bl3 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b3c753 l0bl3 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b3c754 l0bl3 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b3c755 l0bl3 vdd x755 x755b CELLD r1=10000e3 r0=900e3
xl0b3c756 l0bl3 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b3c757 l0bl3 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b3c758 l0bl3 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b3c759 l0bl3 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b3c760 l0bl3 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b3c761 l0bl3 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b3c762 l0bl3 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b3c763 l0bl3 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b3c764 l0bl3 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b3c765 l0bl3 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b3c766 l0bl3 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b3c767 l0bl3 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b3c768 l0bl3 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b3c769 l0bl3 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b3c770 l0bl3 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b3c771 l0bl3 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b3c772 l0bl3 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b3c773 l0bl3 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b3c774 l0bl3 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b3c775 l0bl3 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b3c776 l0bl3 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b3c777 l0bl3 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b3c778 l0bl3 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b3c779 l0bl3 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b3c780 l0bl3 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b3c781 l0bl3 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b3c782 l0bl3 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b3c783 l0bl3 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b4c0 l0bl4 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b4c1 l0bl4 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b4c2 l0bl4 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b4c3 l0bl4 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b4c4 l0bl4 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b4c5 l0bl4 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b4c6 l0bl4 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b4c7 l0bl4 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b4c8 l0bl4 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b4c9 l0bl4 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b4c10 l0bl4 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b4c11 l0bl4 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b4c12 l0bl4 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b4c13 l0bl4 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b4c14 l0bl4 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b4c15 l0bl4 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b4c16 l0bl4 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b4c17 l0bl4 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b4c18 l0bl4 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b4c19 l0bl4 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b4c20 l0bl4 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b4c21 l0bl4 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b4c22 l0bl4 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b4c23 l0bl4 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b4c24 l0bl4 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b4c25 l0bl4 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b4c26 l0bl4 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b4c27 l0bl4 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b4c28 l0bl4 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b4c29 l0bl4 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b4c30 l0bl4 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b4c31 l0bl4 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b4c32 l0bl4 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b4c33 l0bl4 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b4c34 l0bl4 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b4c35 l0bl4 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b4c36 l0bl4 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b4c37 l0bl4 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b4c38 l0bl4 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b4c39 l0bl4 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b4c40 l0bl4 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b4c41 l0bl4 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b4c42 l0bl4 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b4c43 l0bl4 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b4c44 l0bl4 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b4c45 l0bl4 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b4c46 l0bl4 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b4c47 l0bl4 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b4c48 l0bl4 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b4c49 l0bl4 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b4c50 l0bl4 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b4c51 l0bl4 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b4c52 l0bl4 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b4c53 l0bl4 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b4c54 l0bl4 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b4c55 l0bl4 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b4c56 l0bl4 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b4c57 l0bl4 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b4c58 l0bl4 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b4c59 l0bl4 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b4c60 l0bl4 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b4c61 l0bl4 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b4c62 l0bl4 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b4c63 l0bl4 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b4c64 l0bl4 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b4c65 l0bl4 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b4c66 l0bl4 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b4c67 l0bl4 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b4c68 l0bl4 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b4c69 l0bl4 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b4c70 l0bl4 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b4c71 l0bl4 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b4c72 l0bl4 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b4c73 l0bl4 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b4c74 l0bl4 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b4c75 l0bl4 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b4c76 l0bl4 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b4c77 l0bl4 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b4c78 l0bl4 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b4c79 l0bl4 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b4c80 l0bl4 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b4c81 l0bl4 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b4c82 l0bl4 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b4c83 l0bl4 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b4c84 l0bl4 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b4c85 l0bl4 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b4c86 l0bl4 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b4c87 l0bl4 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b4c88 l0bl4 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b4c89 l0bl4 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b4c90 l0bl4 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b4c91 l0bl4 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b4c92 l0bl4 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b4c93 l0bl4 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b4c94 l0bl4 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b4c95 l0bl4 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b4c96 l0bl4 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b4c97 l0bl4 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b4c98 l0bl4 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b4c99 l0bl4 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b4c100 l0bl4 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b4c101 l0bl4 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b4c102 l0bl4 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b4c103 l0bl4 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b4c104 l0bl4 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b4c105 l0bl4 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b4c106 l0bl4 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b4c107 l0bl4 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b4c108 l0bl4 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b4c109 l0bl4 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b4c110 l0bl4 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b4c111 l0bl4 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b4c112 l0bl4 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b4c113 l0bl4 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b4c114 l0bl4 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b4c115 l0bl4 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b4c116 l0bl4 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b4c117 l0bl4 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b4c118 l0bl4 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b4c119 l0bl4 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b4c120 l0bl4 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b4c121 l0bl4 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b4c122 l0bl4 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b4c123 l0bl4 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b4c124 l0bl4 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b4c125 l0bl4 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b4c126 l0bl4 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b4c127 l0bl4 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b4c128 l0bl4 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b4c129 l0bl4 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b4c130 l0bl4 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b4c131 l0bl4 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b4c132 l0bl4 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b4c133 l0bl4 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b4c134 l0bl4 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b4c135 l0bl4 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b4c136 l0bl4 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b4c137 l0bl4 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b4c138 l0bl4 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b4c139 l0bl4 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b4c140 l0bl4 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b4c141 l0bl4 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b4c142 l0bl4 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b4c143 l0bl4 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b4c144 l0bl4 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b4c145 l0bl4 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b4c146 l0bl4 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b4c147 l0bl4 vdd x147 x147b CELLD r1=900e3 r0=10000e3
xl0b4c148 l0bl4 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b4c149 l0bl4 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b4c150 l0bl4 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b4c151 l0bl4 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b4c152 l0bl4 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b4c153 l0bl4 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b4c154 l0bl4 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b4c155 l0bl4 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b4c156 l0bl4 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b4c157 l0bl4 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b4c158 l0bl4 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b4c159 l0bl4 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b4c160 l0bl4 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b4c161 l0bl4 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b4c162 l0bl4 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b4c163 l0bl4 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b4c164 l0bl4 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b4c165 l0bl4 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b4c166 l0bl4 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b4c167 l0bl4 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b4c168 l0bl4 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b4c169 l0bl4 vdd x169 x169b CELLD r1=10000e3 r0=900e3
xl0b4c170 l0bl4 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b4c171 l0bl4 vdd x171 x171b CELLD r1=10000e3 r0=900e3
xl0b4c172 l0bl4 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b4c173 l0bl4 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b4c174 l0bl4 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b4c175 l0bl4 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b4c176 l0bl4 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b4c177 l0bl4 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b4c178 l0bl4 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b4c179 l0bl4 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b4c180 l0bl4 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b4c181 l0bl4 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b4c182 l0bl4 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b4c183 l0bl4 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b4c184 l0bl4 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b4c185 l0bl4 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b4c186 l0bl4 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b4c187 l0bl4 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b4c188 l0bl4 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b4c189 l0bl4 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b4c190 l0bl4 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b4c191 l0bl4 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b4c192 l0bl4 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b4c193 l0bl4 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b4c194 l0bl4 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b4c195 l0bl4 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b4c196 l0bl4 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b4c197 l0bl4 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b4c198 l0bl4 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b4c199 l0bl4 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b4c200 l0bl4 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b4c201 l0bl4 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b4c202 l0bl4 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b4c203 l0bl4 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b4c204 l0bl4 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b4c205 l0bl4 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b4c206 l0bl4 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b4c207 l0bl4 vdd x207 x207b CELLD r1=900e3 r0=10000e3
xl0b4c208 l0bl4 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b4c209 l0bl4 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b4c210 l0bl4 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b4c211 l0bl4 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b4c212 l0bl4 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b4c213 l0bl4 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b4c214 l0bl4 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b4c215 l0bl4 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b4c216 l0bl4 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b4c217 l0bl4 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b4c218 l0bl4 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b4c219 l0bl4 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b4c220 l0bl4 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b4c221 l0bl4 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b4c222 l0bl4 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b4c223 l0bl4 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b4c224 l0bl4 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b4c225 l0bl4 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b4c226 l0bl4 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b4c227 l0bl4 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b4c228 l0bl4 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b4c229 l0bl4 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b4c230 l0bl4 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b4c231 l0bl4 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b4c232 l0bl4 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b4c233 l0bl4 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b4c234 l0bl4 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b4c235 l0bl4 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b4c236 l0bl4 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b4c237 l0bl4 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b4c238 l0bl4 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b4c239 l0bl4 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b4c240 l0bl4 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b4c241 l0bl4 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b4c242 l0bl4 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b4c243 l0bl4 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b4c244 l0bl4 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b4c245 l0bl4 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b4c246 l0bl4 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b4c247 l0bl4 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b4c248 l0bl4 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b4c249 l0bl4 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b4c250 l0bl4 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b4c251 l0bl4 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b4c252 l0bl4 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b4c253 l0bl4 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b4c254 l0bl4 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b4c255 l0bl4 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b4c256 l0bl4 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b4c257 l0bl4 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b4c258 l0bl4 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b4c259 l0bl4 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b4c260 l0bl4 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b4c261 l0bl4 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b4c262 l0bl4 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b4c263 l0bl4 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b4c264 l0bl4 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b4c265 l0bl4 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b4c266 l0bl4 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b4c267 l0bl4 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b4c268 l0bl4 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b4c269 l0bl4 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b4c270 l0bl4 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b4c271 l0bl4 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b4c272 l0bl4 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b4c273 l0bl4 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b4c274 l0bl4 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b4c275 l0bl4 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b4c276 l0bl4 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b4c277 l0bl4 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b4c278 l0bl4 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b4c279 l0bl4 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b4c280 l0bl4 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b4c281 l0bl4 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b4c282 l0bl4 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b4c283 l0bl4 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b4c284 l0bl4 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b4c285 l0bl4 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b4c286 l0bl4 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b4c287 l0bl4 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b4c288 l0bl4 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b4c289 l0bl4 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b4c290 l0bl4 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b4c291 l0bl4 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b4c292 l0bl4 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b4c293 l0bl4 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b4c294 l0bl4 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b4c295 l0bl4 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b4c296 l0bl4 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b4c297 l0bl4 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b4c298 l0bl4 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b4c299 l0bl4 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b4c300 l0bl4 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b4c301 l0bl4 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b4c302 l0bl4 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b4c303 l0bl4 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b4c304 l0bl4 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b4c305 l0bl4 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b4c306 l0bl4 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b4c307 l0bl4 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b4c308 l0bl4 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b4c309 l0bl4 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b4c310 l0bl4 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b4c311 l0bl4 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b4c312 l0bl4 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b4c313 l0bl4 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b4c314 l0bl4 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b4c315 l0bl4 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b4c316 l0bl4 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b4c317 l0bl4 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b4c318 l0bl4 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b4c319 l0bl4 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b4c320 l0bl4 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b4c321 l0bl4 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b4c322 l0bl4 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b4c323 l0bl4 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b4c324 l0bl4 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b4c325 l0bl4 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b4c326 l0bl4 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b4c327 l0bl4 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b4c328 l0bl4 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b4c329 l0bl4 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b4c330 l0bl4 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b4c331 l0bl4 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b4c332 l0bl4 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b4c333 l0bl4 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b4c334 l0bl4 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b4c335 l0bl4 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b4c336 l0bl4 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b4c337 l0bl4 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b4c338 l0bl4 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b4c339 l0bl4 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b4c340 l0bl4 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b4c341 l0bl4 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b4c342 l0bl4 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b4c343 l0bl4 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b4c344 l0bl4 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b4c345 l0bl4 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b4c346 l0bl4 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b4c347 l0bl4 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b4c348 l0bl4 vdd x348 x348b CELLD r1=10000e3 r0=900e3
xl0b4c349 l0bl4 vdd x349 x349b CELLD r1=10000e3 r0=900e3
xl0b4c350 l0bl4 vdd x350 x350b CELLD r1=10000e3 r0=900e3
xl0b4c351 l0bl4 vdd x351 x351b CELLD r1=10000e3 r0=900e3
xl0b4c352 l0bl4 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b4c353 l0bl4 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b4c354 l0bl4 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b4c355 l0bl4 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b4c356 l0bl4 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b4c357 l0bl4 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b4c358 l0bl4 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b4c359 l0bl4 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b4c360 l0bl4 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b4c361 l0bl4 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b4c362 l0bl4 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b4c363 l0bl4 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b4c364 l0bl4 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b4c365 l0bl4 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b4c366 l0bl4 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b4c367 l0bl4 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b4c368 l0bl4 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b4c369 l0bl4 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b4c370 l0bl4 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b4c371 l0bl4 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b4c372 l0bl4 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b4c373 l0bl4 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b4c374 l0bl4 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b4c375 l0bl4 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b4c376 l0bl4 vdd x376 x376b CELLD r1=10000e3 r0=900e3
xl0b4c377 l0bl4 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b4c378 l0bl4 vdd x378 x378b CELLD r1=10000e3 r0=900e3
xl0b4c379 l0bl4 vdd x379 x379b CELLD r1=10000e3 r0=900e3
xl0b4c380 l0bl4 vdd x380 x380b CELLD r1=10000e3 r0=900e3
xl0b4c381 l0bl4 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b4c382 l0bl4 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b4c383 l0bl4 vdd x383 x383b CELLD r1=10000e3 r0=900e3
xl0b4c384 l0bl4 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b4c385 l0bl4 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b4c386 l0bl4 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b4c387 l0bl4 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b4c388 l0bl4 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b4c389 l0bl4 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b4c390 l0bl4 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b4c391 l0bl4 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b4c392 l0bl4 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b4c393 l0bl4 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b4c394 l0bl4 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b4c395 l0bl4 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b4c396 l0bl4 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b4c397 l0bl4 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b4c398 l0bl4 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b4c399 l0bl4 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b4c400 l0bl4 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b4c401 l0bl4 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b4c402 l0bl4 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b4c403 l0bl4 vdd x403 x403b CELLD r1=10000e3 r0=900e3
xl0b4c404 l0bl4 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b4c405 l0bl4 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b4c406 l0bl4 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b4c407 l0bl4 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b4c408 l0bl4 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b4c409 l0bl4 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b4c410 l0bl4 vdd x410 x410b CELLD r1=10000e3 r0=900e3
xl0b4c411 l0bl4 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b4c412 l0bl4 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b4c413 l0bl4 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b4c414 l0bl4 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b4c415 l0bl4 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b4c416 l0bl4 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b4c417 l0bl4 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b4c418 l0bl4 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b4c419 l0bl4 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b4c420 l0bl4 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b4c421 l0bl4 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b4c422 l0bl4 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b4c423 l0bl4 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b4c424 l0bl4 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b4c425 l0bl4 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b4c426 l0bl4 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b4c427 l0bl4 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b4c428 l0bl4 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b4c429 l0bl4 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b4c430 l0bl4 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b4c431 l0bl4 vdd x431 x431b CELLD r1=10000e3 r0=900e3
xl0b4c432 l0bl4 vdd x432 x432b CELLD r1=10000e3 r0=900e3
xl0b4c433 l0bl4 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b4c434 l0bl4 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b4c435 l0bl4 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b4c436 l0bl4 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b4c437 l0bl4 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b4c438 l0bl4 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b4c439 l0bl4 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b4c440 l0bl4 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b4c441 l0bl4 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b4c442 l0bl4 vdd x442 x442b CELLD r1=900e3 r0=10000e3
xl0b4c443 l0bl4 vdd x443 x443b CELLD r1=900e3 r0=10000e3
xl0b4c444 l0bl4 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b4c445 l0bl4 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b4c446 l0bl4 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b4c447 l0bl4 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b4c448 l0bl4 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b4c449 l0bl4 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b4c450 l0bl4 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b4c451 l0bl4 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b4c452 l0bl4 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b4c453 l0bl4 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b4c454 l0bl4 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b4c455 l0bl4 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b4c456 l0bl4 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b4c457 l0bl4 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b4c458 l0bl4 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b4c459 l0bl4 vdd x459 x459b CELLD r1=10000e3 r0=900e3
xl0b4c460 l0bl4 vdd x460 x460b CELLD r1=10000e3 r0=900e3
xl0b4c461 l0bl4 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b4c462 l0bl4 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b4c463 l0bl4 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b4c464 l0bl4 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b4c465 l0bl4 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b4c466 l0bl4 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b4c467 l0bl4 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b4c468 l0bl4 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b4c469 l0bl4 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b4c470 l0bl4 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b4c471 l0bl4 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b4c472 l0bl4 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b4c473 l0bl4 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b4c474 l0bl4 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b4c475 l0bl4 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b4c476 l0bl4 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b4c477 l0bl4 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b4c478 l0bl4 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b4c479 l0bl4 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b4c480 l0bl4 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b4c481 l0bl4 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b4c482 l0bl4 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b4c483 l0bl4 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b4c484 l0bl4 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b4c485 l0bl4 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b4c486 l0bl4 vdd x486 x486b CELLD r1=10000e3 r0=900e3
xl0b4c487 l0bl4 vdd x487 x487b CELLD r1=10000e3 r0=900e3
xl0b4c488 l0bl4 vdd x488 x488b CELLD r1=10000e3 r0=900e3
xl0b4c489 l0bl4 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b4c490 l0bl4 vdd x490 x490b CELLD r1=10000e3 r0=900e3
xl0b4c491 l0bl4 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b4c492 l0bl4 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b4c493 l0bl4 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b4c494 l0bl4 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b4c495 l0bl4 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b4c496 l0bl4 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b4c497 l0bl4 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b4c498 l0bl4 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b4c499 l0bl4 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b4c500 l0bl4 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b4c501 l0bl4 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b4c502 l0bl4 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b4c503 l0bl4 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b4c504 l0bl4 vdd x504 x504b CELLD r1=10000e3 r0=900e3
xl0b4c505 l0bl4 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b4c506 l0bl4 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b4c507 l0bl4 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b4c508 l0bl4 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b4c509 l0bl4 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b4c510 l0bl4 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b4c511 l0bl4 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b4c512 l0bl4 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b4c513 l0bl4 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b4c514 l0bl4 vdd x514 x514b CELLD r1=10000e3 r0=900e3
xl0b4c515 l0bl4 vdd x515 x515b CELLD r1=10000e3 r0=900e3
xl0b4c516 l0bl4 vdd x516 x516b CELLD r1=10000e3 r0=900e3
xl0b4c517 l0bl4 vdd x517 x517b CELLD r1=10000e3 r0=900e3
xl0b4c518 l0bl4 vdd x518 x518b CELLD r1=10000e3 r0=900e3
xl0b4c519 l0bl4 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b4c520 l0bl4 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b4c521 l0bl4 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b4c522 l0bl4 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b4c523 l0bl4 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b4c524 l0bl4 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b4c525 l0bl4 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b4c526 l0bl4 vdd x526 x526b CELLD r1=900e3 r0=10000e3
xl0b4c527 l0bl4 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b4c528 l0bl4 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b4c529 l0bl4 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b4c530 l0bl4 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b4c531 l0bl4 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b4c532 l0bl4 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b4c533 l0bl4 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b4c534 l0bl4 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b4c535 l0bl4 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b4c536 l0bl4 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b4c537 l0bl4 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b4c538 l0bl4 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b4c539 l0bl4 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b4c540 l0bl4 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b4c541 l0bl4 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b4c542 l0bl4 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b4c543 l0bl4 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b4c544 l0bl4 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b4c545 l0bl4 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b4c546 l0bl4 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b4c547 l0bl4 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b4c548 l0bl4 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b4c549 l0bl4 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b4c550 l0bl4 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b4c551 l0bl4 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b4c552 l0bl4 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b4c553 l0bl4 vdd x553 x553b CELLD r1=900e3 r0=10000e3
xl0b4c554 l0bl4 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b4c555 l0bl4 vdd x555 x555b CELLD r1=900e3 r0=10000e3
xl0b4c556 l0bl4 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b4c557 l0bl4 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b4c558 l0bl4 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b4c559 l0bl4 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b4c560 l0bl4 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b4c561 l0bl4 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b4c562 l0bl4 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b4c563 l0bl4 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b4c564 l0bl4 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b4c565 l0bl4 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b4c566 l0bl4 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b4c567 l0bl4 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b4c568 l0bl4 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b4c569 l0bl4 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b4c570 l0bl4 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b4c571 l0bl4 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b4c572 l0bl4 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b4c573 l0bl4 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b4c574 l0bl4 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b4c575 l0bl4 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b4c576 l0bl4 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b4c577 l0bl4 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b4c578 l0bl4 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b4c579 l0bl4 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b4c580 l0bl4 vdd x580 x580b CELLD r1=900e3 r0=10000e3
xl0b4c581 l0bl4 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b4c582 l0bl4 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b4c583 l0bl4 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b4c584 l0bl4 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b4c585 l0bl4 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b4c586 l0bl4 vdd x586 x586b CELLD r1=10000e3 r0=900e3
xl0b4c587 l0bl4 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b4c588 l0bl4 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b4c589 l0bl4 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b4c590 l0bl4 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b4c591 l0bl4 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b4c592 l0bl4 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b4c593 l0bl4 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b4c594 l0bl4 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b4c595 l0bl4 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b4c596 l0bl4 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b4c597 l0bl4 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b4c598 l0bl4 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b4c599 l0bl4 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b4c600 l0bl4 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b4c601 l0bl4 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b4c602 l0bl4 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b4c603 l0bl4 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b4c604 l0bl4 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b4c605 l0bl4 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b4c606 l0bl4 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b4c607 l0bl4 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b4c608 l0bl4 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b4c609 l0bl4 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b4c610 l0bl4 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b4c611 l0bl4 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b4c612 l0bl4 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b4c613 l0bl4 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b4c614 l0bl4 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b4c615 l0bl4 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b4c616 l0bl4 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b4c617 l0bl4 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b4c618 l0bl4 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b4c619 l0bl4 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b4c620 l0bl4 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b4c621 l0bl4 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b4c622 l0bl4 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b4c623 l0bl4 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b4c624 l0bl4 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b4c625 l0bl4 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b4c626 l0bl4 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b4c627 l0bl4 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b4c628 l0bl4 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b4c629 l0bl4 vdd x629 x629b CELLD r1=900e3 r0=10000e3
xl0b4c630 l0bl4 vdd x630 x630b CELLD r1=900e3 r0=10000e3
xl0b4c631 l0bl4 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b4c632 l0bl4 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b4c633 l0bl4 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b4c634 l0bl4 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b4c635 l0bl4 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b4c636 l0bl4 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b4c637 l0bl4 vdd x637 x637b CELLD r1=10000e3 r0=900e3
xl0b4c638 l0bl4 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b4c639 l0bl4 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b4c640 l0bl4 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b4c641 l0bl4 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b4c642 l0bl4 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b4c643 l0bl4 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b4c644 l0bl4 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b4c645 l0bl4 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b4c646 l0bl4 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b4c647 l0bl4 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b4c648 l0bl4 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b4c649 l0bl4 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b4c650 l0bl4 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b4c651 l0bl4 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b4c652 l0bl4 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b4c653 l0bl4 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b4c654 l0bl4 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b4c655 l0bl4 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b4c656 l0bl4 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b4c657 l0bl4 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b4c658 l0bl4 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b4c659 l0bl4 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b4c660 l0bl4 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b4c661 l0bl4 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b4c662 l0bl4 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b4c663 l0bl4 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b4c664 l0bl4 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b4c665 l0bl4 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b4c666 l0bl4 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b4c667 l0bl4 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b4c668 l0bl4 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b4c669 l0bl4 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b4c670 l0bl4 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b4c671 l0bl4 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b4c672 l0bl4 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b4c673 l0bl4 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b4c674 l0bl4 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b4c675 l0bl4 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b4c676 l0bl4 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b4c677 l0bl4 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b4c678 l0bl4 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b4c679 l0bl4 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b4c680 l0bl4 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b4c681 l0bl4 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b4c682 l0bl4 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b4c683 l0bl4 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b4c684 l0bl4 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b4c685 l0bl4 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b4c686 l0bl4 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b4c687 l0bl4 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b4c688 l0bl4 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b4c689 l0bl4 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b4c690 l0bl4 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b4c691 l0bl4 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b4c692 l0bl4 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b4c693 l0bl4 vdd x693 x693b CELLD r1=10000e3 r0=900e3
xl0b4c694 l0bl4 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b4c695 l0bl4 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b4c696 l0bl4 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b4c697 l0bl4 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b4c698 l0bl4 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b4c699 l0bl4 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b4c700 l0bl4 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b4c701 l0bl4 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b4c702 l0bl4 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b4c703 l0bl4 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b4c704 l0bl4 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b4c705 l0bl4 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b4c706 l0bl4 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b4c707 l0bl4 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b4c708 l0bl4 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b4c709 l0bl4 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b4c710 l0bl4 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b4c711 l0bl4 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b4c712 l0bl4 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b4c713 l0bl4 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b4c714 l0bl4 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b4c715 l0bl4 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b4c716 l0bl4 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b4c717 l0bl4 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b4c718 l0bl4 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b4c719 l0bl4 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b4c720 l0bl4 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b4c721 l0bl4 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b4c722 l0bl4 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b4c723 l0bl4 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b4c724 l0bl4 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b4c725 l0bl4 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b4c726 l0bl4 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b4c727 l0bl4 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b4c728 l0bl4 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b4c729 l0bl4 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b4c730 l0bl4 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b4c731 l0bl4 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b4c732 l0bl4 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b4c733 l0bl4 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b4c734 l0bl4 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b4c735 l0bl4 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b4c736 l0bl4 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b4c737 l0bl4 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b4c738 l0bl4 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b4c739 l0bl4 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b4c740 l0bl4 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b4c741 l0bl4 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b4c742 l0bl4 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b4c743 l0bl4 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b4c744 l0bl4 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b4c745 l0bl4 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b4c746 l0bl4 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b4c747 l0bl4 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b4c748 l0bl4 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b4c749 l0bl4 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b4c750 l0bl4 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b4c751 l0bl4 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b4c752 l0bl4 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b4c753 l0bl4 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b4c754 l0bl4 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b4c755 l0bl4 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b4c756 l0bl4 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b4c757 l0bl4 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b4c758 l0bl4 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b4c759 l0bl4 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b4c760 l0bl4 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b4c761 l0bl4 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b4c762 l0bl4 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b4c763 l0bl4 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b4c764 l0bl4 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b4c765 l0bl4 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b4c766 l0bl4 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b4c767 l0bl4 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b4c768 l0bl4 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b4c769 l0bl4 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b4c770 l0bl4 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b4c771 l0bl4 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b4c772 l0bl4 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b4c773 l0bl4 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b4c774 l0bl4 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b4c775 l0bl4 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b4c776 l0bl4 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b4c777 l0bl4 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b4c778 l0bl4 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b4c779 l0bl4 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b4c780 l0bl4 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b4c781 l0bl4 vdd x781 x781b CELLD r1=10000e3 r0=900e3
xl0b4c782 l0bl4 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b4c783 l0bl4 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b5c0 l0bl5 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b5c1 l0bl5 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b5c2 l0bl5 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b5c3 l0bl5 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b5c4 l0bl5 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b5c5 l0bl5 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b5c6 l0bl5 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b5c7 l0bl5 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b5c8 l0bl5 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b5c9 l0bl5 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b5c10 l0bl5 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b5c11 l0bl5 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b5c12 l0bl5 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b5c13 l0bl5 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b5c14 l0bl5 vdd x14 x14b CELLD r1=10000e3 r0=900e3
xl0b5c15 l0bl5 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b5c16 l0bl5 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b5c17 l0bl5 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b5c18 l0bl5 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b5c19 l0bl5 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b5c20 l0bl5 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b5c21 l0bl5 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b5c22 l0bl5 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b5c23 l0bl5 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b5c24 l0bl5 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b5c25 l0bl5 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b5c26 l0bl5 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b5c27 l0bl5 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b5c28 l0bl5 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b5c29 l0bl5 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b5c30 l0bl5 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b5c31 l0bl5 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b5c32 l0bl5 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b5c33 l0bl5 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b5c34 l0bl5 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b5c35 l0bl5 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b5c36 l0bl5 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b5c37 l0bl5 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b5c38 l0bl5 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b5c39 l0bl5 vdd x39 x39b CELLD r1=10000e3 r0=900e3
xl0b5c40 l0bl5 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b5c41 l0bl5 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b5c42 l0bl5 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b5c43 l0bl5 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b5c44 l0bl5 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b5c45 l0bl5 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b5c46 l0bl5 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b5c47 l0bl5 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b5c48 l0bl5 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b5c49 l0bl5 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b5c50 l0bl5 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b5c51 l0bl5 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b5c52 l0bl5 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b5c53 l0bl5 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b5c54 l0bl5 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b5c55 l0bl5 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b5c56 l0bl5 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b5c57 l0bl5 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b5c58 l0bl5 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b5c59 l0bl5 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b5c60 l0bl5 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b5c61 l0bl5 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b5c62 l0bl5 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b5c63 l0bl5 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b5c64 l0bl5 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b5c65 l0bl5 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b5c66 l0bl5 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b5c67 l0bl5 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b5c68 l0bl5 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b5c69 l0bl5 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b5c70 l0bl5 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b5c71 l0bl5 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b5c72 l0bl5 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b5c73 l0bl5 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b5c74 l0bl5 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b5c75 l0bl5 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b5c76 l0bl5 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b5c77 l0bl5 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b5c78 l0bl5 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b5c79 l0bl5 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b5c80 l0bl5 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b5c81 l0bl5 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b5c82 l0bl5 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b5c83 l0bl5 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b5c84 l0bl5 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b5c85 l0bl5 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b5c86 l0bl5 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b5c87 l0bl5 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b5c88 l0bl5 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b5c89 l0bl5 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b5c90 l0bl5 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b5c91 l0bl5 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b5c92 l0bl5 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b5c93 l0bl5 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b5c94 l0bl5 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b5c95 l0bl5 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b5c96 l0bl5 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b5c97 l0bl5 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b5c98 l0bl5 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b5c99 l0bl5 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b5c100 l0bl5 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b5c101 l0bl5 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b5c102 l0bl5 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b5c103 l0bl5 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b5c104 l0bl5 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b5c105 l0bl5 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b5c106 l0bl5 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b5c107 l0bl5 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b5c108 l0bl5 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b5c109 l0bl5 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b5c110 l0bl5 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b5c111 l0bl5 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b5c112 l0bl5 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b5c113 l0bl5 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b5c114 l0bl5 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b5c115 l0bl5 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b5c116 l0bl5 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b5c117 l0bl5 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b5c118 l0bl5 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b5c119 l0bl5 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b5c120 l0bl5 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b5c121 l0bl5 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b5c122 l0bl5 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b5c123 l0bl5 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b5c124 l0bl5 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b5c125 l0bl5 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b5c126 l0bl5 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b5c127 l0bl5 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b5c128 l0bl5 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b5c129 l0bl5 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b5c130 l0bl5 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b5c131 l0bl5 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b5c132 l0bl5 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b5c133 l0bl5 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b5c134 l0bl5 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b5c135 l0bl5 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b5c136 l0bl5 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b5c137 l0bl5 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b5c138 l0bl5 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b5c139 l0bl5 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b5c140 l0bl5 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b5c141 l0bl5 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b5c142 l0bl5 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b5c143 l0bl5 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b5c144 l0bl5 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b5c145 l0bl5 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b5c146 l0bl5 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b5c147 l0bl5 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b5c148 l0bl5 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b5c149 l0bl5 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b5c150 l0bl5 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b5c151 l0bl5 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b5c152 l0bl5 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b5c153 l0bl5 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b5c154 l0bl5 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b5c155 l0bl5 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b5c156 l0bl5 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b5c157 l0bl5 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b5c158 l0bl5 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b5c159 l0bl5 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b5c160 l0bl5 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b5c161 l0bl5 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b5c162 l0bl5 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b5c163 l0bl5 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b5c164 l0bl5 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b5c165 l0bl5 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b5c166 l0bl5 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b5c167 l0bl5 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b5c168 l0bl5 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b5c169 l0bl5 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b5c170 l0bl5 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b5c171 l0bl5 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b5c172 l0bl5 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b5c173 l0bl5 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b5c174 l0bl5 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b5c175 l0bl5 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b5c176 l0bl5 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b5c177 l0bl5 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b5c178 l0bl5 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b5c179 l0bl5 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b5c180 l0bl5 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b5c181 l0bl5 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b5c182 l0bl5 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b5c183 l0bl5 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b5c184 l0bl5 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b5c185 l0bl5 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b5c186 l0bl5 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b5c187 l0bl5 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b5c188 l0bl5 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b5c189 l0bl5 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b5c190 l0bl5 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b5c191 l0bl5 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b5c192 l0bl5 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b5c193 l0bl5 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b5c194 l0bl5 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b5c195 l0bl5 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b5c196 l0bl5 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b5c197 l0bl5 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b5c198 l0bl5 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b5c199 l0bl5 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b5c200 l0bl5 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b5c201 l0bl5 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b5c202 l0bl5 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b5c203 l0bl5 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b5c204 l0bl5 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b5c205 l0bl5 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b5c206 l0bl5 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b5c207 l0bl5 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b5c208 l0bl5 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b5c209 l0bl5 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b5c210 l0bl5 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b5c211 l0bl5 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b5c212 l0bl5 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b5c213 l0bl5 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b5c214 l0bl5 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b5c215 l0bl5 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b5c216 l0bl5 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b5c217 l0bl5 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b5c218 l0bl5 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b5c219 l0bl5 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b5c220 l0bl5 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b5c221 l0bl5 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b5c222 l0bl5 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b5c223 l0bl5 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b5c224 l0bl5 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b5c225 l0bl5 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b5c226 l0bl5 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b5c227 l0bl5 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b5c228 l0bl5 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b5c229 l0bl5 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b5c230 l0bl5 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b5c231 l0bl5 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b5c232 l0bl5 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b5c233 l0bl5 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b5c234 l0bl5 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b5c235 l0bl5 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b5c236 l0bl5 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b5c237 l0bl5 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b5c238 l0bl5 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b5c239 l0bl5 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b5c240 l0bl5 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b5c241 l0bl5 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b5c242 l0bl5 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b5c243 l0bl5 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b5c244 l0bl5 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b5c245 l0bl5 vdd x245 x245b CELLD r1=900e3 r0=10000e3
xl0b5c246 l0bl5 vdd x246 x246b CELLD r1=900e3 r0=10000e3
xl0b5c247 l0bl5 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b5c248 l0bl5 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b5c249 l0bl5 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b5c250 l0bl5 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b5c251 l0bl5 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b5c252 l0bl5 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b5c253 l0bl5 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b5c254 l0bl5 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b5c255 l0bl5 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b5c256 l0bl5 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b5c257 l0bl5 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b5c258 l0bl5 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b5c259 l0bl5 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b5c260 l0bl5 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b5c261 l0bl5 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b5c262 l0bl5 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b5c263 l0bl5 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b5c264 l0bl5 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b5c265 l0bl5 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b5c266 l0bl5 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b5c267 l0bl5 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b5c268 l0bl5 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b5c269 l0bl5 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b5c270 l0bl5 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b5c271 l0bl5 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b5c272 l0bl5 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b5c273 l0bl5 vdd x273 x273b CELLD r1=900e3 r0=10000e3
xl0b5c274 l0bl5 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b5c275 l0bl5 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b5c276 l0bl5 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b5c277 l0bl5 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b5c278 l0bl5 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b5c279 l0bl5 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b5c280 l0bl5 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b5c281 l0bl5 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b5c282 l0bl5 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b5c283 l0bl5 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b5c284 l0bl5 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b5c285 l0bl5 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b5c286 l0bl5 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b5c287 l0bl5 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b5c288 l0bl5 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b5c289 l0bl5 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b5c290 l0bl5 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b5c291 l0bl5 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b5c292 l0bl5 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b5c293 l0bl5 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b5c294 l0bl5 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b5c295 l0bl5 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b5c296 l0bl5 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b5c297 l0bl5 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b5c298 l0bl5 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b5c299 l0bl5 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b5c300 l0bl5 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b5c301 l0bl5 vdd x301 x301b CELLD r1=900e3 r0=10000e3
xl0b5c302 l0bl5 vdd x302 x302b CELLD r1=900e3 r0=10000e3
xl0b5c303 l0bl5 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b5c304 l0bl5 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b5c305 l0bl5 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b5c306 l0bl5 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b5c307 l0bl5 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b5c308 l0bl5 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b5c309 l0bl5 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b5c310 l0bl5 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b5c311 l0bl5 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b5c312 l0bl5 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b5c313 l0bl5 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b5c314 l0bl5 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b5c315 l0bl5 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b5c316 l0bl5 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b5c317 l0bl5 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b5c318 l0bl5 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b5c319 l0bl5 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b5c320 l0bl5 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b5c321 l0bl5 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b5c322 l0bl5 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b5c323 l0bl5 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b5c324 l0bl5 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b5c325 l0bl5 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b5c326 l0bl5 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b5c327 l0bl5 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b5c328 l0bl5 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b5c329 l0bl5 vdd x329 x329b CELLD r1=900e3 r0=10000e3
xl0b5c330 l0bl5 vdd x330 x330b CELLD r1=900e3 r0=10000e3
xl0b5c331 l0bl5 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b5c332 l0bl5 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b5c333 l0bl5 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b5c334 l0bl5 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b5c335 l0bl5 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b5c336 l0bl5 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b5c337 l0bl5 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b5c338 l0bl5 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b5c339 l0bl5 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b5c340 l0bl5 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b5c341 l0bl5 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b5c342 l0bl5 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b5c343 l0bl5 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b5c344 l0bl5 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b5c345 l0bl5 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b5c346 l0bl5 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b5c347 l0bl5 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b5c348 l0bl5 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b5c349 l0bl5 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b5c350 l0bl5 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b5c351 l0bl5 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b5c352 l0bl5 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b5c353 l0bl5 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b5c354 l0bl5 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b5c355 l0bl5 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b5c356 l0bl5 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b5c357 l0bl5 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b5c358 l0bl5 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b5c359 l0bl5 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b5c360 l0bl5 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b5c361 l0bl5 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b5c362 l0bl5 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b5c363 l0bl5 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b5c364 l0bl5 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b5c365 l0bl5 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b5c366 l0bl5 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b5c367 l0bl5 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b5c368 l0bl5 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b5c369 l0bl5 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b5c370 l0bl5 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b5c371 l0bl5 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b5c372 l0bl5 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b5c373 l0bl5 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b5c374 l0bl5 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b5c375 l0bl5 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b5c376 l0bl5 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b5c377 l0bl5 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b5c378 l0bl5 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b5c379 l0bl5 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b5c380 l0bl5 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b5c381 l0bl5 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b5c382 l0bl5 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b5c383 l0bl5 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b5c384 l0bl5 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b5c385 l0bl5 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b5c386 l0bl5 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b5c387 l0bl5 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b5c388 l0bl5 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b5c389 l0bl5 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b5c390 l0bl5 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b5c391 l0bl5 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b5c392 l0bl5 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b5c393 l0bl5 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b5c394 l0bl5 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b5c395 l0bl5 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b5c396 l0bl5 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b5c397 l0bl5 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b5c398 l0bl5 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b5c399 l0bl5 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b5c400 l0bl5 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b5c401 l0bl5 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b5c402 l0bl5 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b5c403 l0bl5 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b5c404 l0bl5 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b5c405 l0bl5 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b5c406 l0bl5 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b5c407 l0bl5 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b5c408 l0bl5 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b5c409 l0bl5 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b5c410 l0bl5 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b5c411 l0bl5 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b5c412 l0bl5 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b5c413 l0bl5 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b5c414 l0bl5 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b5c415 l0bl5 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b5c416 l0bl5 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b5c417 l0bl5 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b5c418 l0bl5 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b5c419 l0bl5 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b5c420 l0bl5 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b5c421 l0bl5 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b5c422 l0bl5 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b5c423 l0bl5 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b5c424 l0bl5 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b5c425 l0bl5 vdd x425 x425b CELLD r1=900e3 r0=10000e3
xl0b5c426 l0bl5 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b5c427 l0bl5 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b5c428 l0bl5 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b5c429 l0bl5 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b5c430 l0bl5 vdd x430 x430b CELLD r1=10000e3 r0=900e3
xl0b5c431 l0bl5 vdd x431 x431b CELLD r1=10000e3 r0=900e3
xl0b5c432 l0bl5 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b5c433 l0bl5 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b5c434 l0bl5 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b5c435 l0bl5 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b5c436 l0bl5 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b5c437 l0bl5 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b5c438 l0bl5 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b5c439 l0bl5 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b5c440 l0bl5 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b5c441 l0bl5 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b5c442 l0bl5 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b5c443 l0bl5 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b5c444 l0bl5 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b5c445 l0bl5 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b5c446 l0bl5 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b5c447 l0bl5 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b5c448 l0bl5 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b5c449 l0bl5 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b5c450 l0bl5 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b5c451 l0bl5 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b5c452 l0bl5 vdd x452 x452b CELLD r1=900e3 r0=10000e3
xl0b5c453 l0bl5 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b5c454 l0bl5 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b5c455 l0bl5 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b5c456 l0bl5 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b5c457 l0bl5 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b5c458 l0bl5 vdd x458 x458b CELLD r1=10000e3 r0=900e3
xl0b5c459 l0bl5 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b5c460 l0bl5 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b5c461 l0bl5 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b5c462 l0bl5 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b5c463 l0bl5 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b5c464 l0bl5 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b5c465 l0bl5 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b5c466 l0bl5 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b5c467 l0bl5 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b5c468 l0bl5 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b5c469 l0bl5 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b5c470 l0bl5 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b5c471 l0bl5 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b5c472 l0bl5 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b5c473 l0bl5 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b5c474 l0bl5 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b5c475 l0bl5 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b5c476 l0bl5 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b5c477 l0bl5 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b5c478 l0bl5 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b5c479 l0bl5 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b5c480 l0bl5 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b5c481 l0bl5 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b5c482 l0bl5 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b5c483 l0bl5 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b5c484 l0bl5 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b5c485 l0bl5 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b5c486 l0bl5 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b5c487 l0bl5 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b5c488 l0bl5 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b5c489 l0bl5 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b5c490 l0bl5 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b5c491 l0bl5 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b5c492 l0bl5 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b5c493 l0bl5 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b5c494 l0bl5 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b5c495 l0bl5 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b5c496 l0bl5 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b5c497 l0bl5 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b5c498 l0bl5 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b5c499 l0bl5 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b5c500 l0bl5 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b5c501 l0bl5 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b5c502 l0bl5 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b5c503 l0bl5 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b5c504 l0bl5 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b5c505 l0bl5 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b5c506 l0bl5 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b5c507 l0bl5 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b5c508 l0bl5 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b5c509 l0bl5 vdd x509 x509b CELLD r1=900e3 r0=10000e3
xl0b5c510 l0bl5 vdd x510 x510b CELLD r1=900e3 r0=10000e3
xl0b5c511 l0bl5 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b5c512 l0bl5 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b5c513 l0bl5 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b5c514 l0bl5 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b5c515 l0bl5 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b5c516 l0bl5 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b5c517 l0bl5 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b5c518 l0bl5 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b5c519 l0bl5 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b5c520 l0bl5 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b5c521 l0bl5 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b5c522 l0bl5 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b5c523 l0bl5 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b5c524 l0bl5 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b5c525 l0bl5 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b5c526 l0bl5 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b5c527 l0bl5 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b5c528 l0bl5 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b5c529 l0bl5 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b5c530 l0bl5 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b5c531 l0bl5 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b5c532 l0bl5 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b5c533 l0bl5 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b5c534 l0bl5 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b5c535 l0bl5 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b5c536 l0bl5 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b5c537 l0bl5 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b5c538 l0bl5 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b5c539 l0bl5 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b5c540 l0bl5 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b5c541 l0bl5 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b5c542 l0bl5 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b5c543 l0bl5 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b5c544 l0bl5 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b5c545 l0bl5 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b5c546 l0bl5 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b5c547 l0bl5 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b5c548 l0bl5 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b5c549 l0bl5 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b5c550 l0bl5 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b5c551 l0bl5 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b5c552 l0bl5 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b5c553 l0bl5 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b5c554 l0bl5 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b5c555 l0bl5 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b5c556 l0bl5 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b5c557 l0bl5 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b5c558 l0bl5 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b5c559 l0bl5 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b5c560 l0bl5 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b5c561 l0bl5 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b5c562 l0bl5 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b5c563 l0bl5 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b5c564 l0bl5 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b5c565 l0bl5 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b5c566 l0bl5 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b5c567 l0bl5 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b5c568 l0bl5 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b5c569 l0bl5 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b5c570 l0bl5 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b5c571 l0bl5 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b5c572 l0bl5 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b5c573 l0bl5 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b5c574 l0bl5 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b5c575 l0bl5 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b5c576 l0bl5 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b5c577 l0bl5 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b5c578 l0bl5 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b5c579 l0bl5 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b5c580 l0bl5 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b5c581 l0bl5 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b5c582 l0bl5 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b5c583 l0bl5 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b5c584 l0bl5 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b5c585 l0bl5 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b5c586 l0bl5 vdd x586 x586b CELLD r1=10000e3 r0=900e3
xl0b5c587 l0bl5 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b5c588 l0bl5 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b5c589 l0bl5 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b5c590 l0bl5 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b5c591 l0bl5 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b5c592 l0bl5 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b5c593 l0bl5 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b5c594 l0bl5 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b5c595 l0bl5 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b5c596 l0bl5 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b5c597 l0bl5 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b5c598 l0bl5 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b5c599 l0bl5 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b5c600 l0bl5 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b5c601 l0bl5 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b5c602 l0bl5 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b5c603 l0bl5 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b5c604 l0bl5 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b5c605 l0bl5 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b5c606 l0bl5 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b5c607 l0bl5 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b5c608 l0bl5 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b5c609 l0bl5 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b5c610 l0bl5 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b5c611 l0bl5 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b5c612 l0bl5 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b5c613 l0bl5 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b5c614 l0bl5 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b5c615 l0bl5 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b5c616 l0bl5 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b5c617 l0bl5 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b5c618 l0bl5 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b5c619 l0bl5 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b5c620 l0bl5 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b5c621 l0bl5 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b5c622 l0bl5 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b5c623 l0bl5 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b5c624 l0bl5 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b5c625 l0bl5 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b5c626 l0bl5 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b5c627 l0bl5 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b5c628 l0bl5 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b5c629 l0bl5 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b5c630 l0bl5 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b5c631 l0bl5 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b5c632 l0bl5 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b5c633 l0bl5 vdd x633 x633b CELLD r1=10000e3 r0=900e3
xl0b5c634 l0bl5 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b5c635 l0bl5 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b5c636 l0bl5 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b5c637 l0bl5 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b5c638 l0bl5 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b5c639 l0bl5 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b5c640 l0bl5 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b5c641 l0bl5 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b5c642 l0bl5 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b5c643 l0bl5 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b5c644 l0bl5 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b5c645 l0bl5 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b5c646 l0bl5 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b5c647 l0bl5 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b5c648 l0bl5 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b5c649 l0bl5 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b5c650 l0bl5 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b5c651 l0bl5 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b5c652 l0bl5 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b5c653 l0bl5 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b5c654 l0bl5 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b5c655 l0bl5 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b5c656 l0bl5 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b5c657 l0bl5 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b5c658 l0bl5 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b5c659 l0bl5 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b5c660 l0bl5 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b5c661 l0bl5 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b5c662 l0bl5 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b5c663 l0bl5 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b5c664 l0bl5 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b5c665 l0bl5 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b5c666 l0bl5 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b5c667 l0bl5 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b5c668 l0bl5 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b5c669 l0bl5 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b5c670 l0bl5 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b5c671 l0bl5 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b5c672 l0bl5 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b5c673 l0bl5 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b5c674 l0bl5 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b5c675 l0bl5 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b5c676 l0bl5 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b5c677 l0bl5 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b5c678 l0bl5 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b5c679 l0bl5 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b5c680 l0bl5 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b5c681 l0bl5 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b5c682 l0bl5 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b5c683 l0bl5 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b5c684 l0bl5 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b5c685 l0bl5 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b5c686 l0bl5 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b5c687 l0bl5 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b5c688 l0bl5 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b5c689 l0bl5 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b5c690 l0bl5 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b5c691 l0bl5 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b5c692 l0bl5 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b5c693 l0bl5 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b5c694 l0bl5 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b5c695 l0bl5 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b5c696 l0bl5 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b5c697 l0bl5 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b5c698 l0bl5 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b5c699 l0bl5 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b5c700 l0bl5 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b5c701 l0bl5 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b5c702 l0bl5 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b5c703 l0bl5 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b5c704 l0bl5 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b5c705 l0bl5 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b5c706 l0bl5 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b5c707 l0bl5 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b5c708 l0bl5 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b5c709 l0bl5 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b5c710 l0bl5 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b5c711 l0bl5 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b5c712 l0bl5 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b5c713 l0bl5 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b5c714 l0bl5 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b5c715 l0bl5 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b5c716 l0bl5 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b5c717 l0bl5 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b5c718 l0bl5 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b5c719 l0bl5 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b5c720 l0bl5 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b5c721 l0bl5 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b5c722 l0bl5 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b5c723 l0bl5 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b5c724 l0bl5 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b5c725 l0bl5 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b5c726 l0bl5 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b5c727 l0bl5 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b5c728 l0bl5 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b5c729 l0bl5 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b5c730 l0bl5 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b5c731 l0bl5 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b5c732 l0bl5 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b5c733 l0bl5 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b5c734 l0bl5 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b5c735 l0bl5 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b5c736 l0bl5 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b5c737 l0bl5 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b5c738 l0bl5 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b5c739 l0bl5 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b5c740 l0bl5 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b5c741 l0bl5 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b5c742 l0bl5 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b5c743 l0bl5 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b5c744 l0bl5 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b5c745 l0bl5 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b5c746 l0bl5 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b5c747 l0bl5 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b5c748 l0bl5 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b5c749 l0bl5 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b5c750 l0bl5 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b5c751 l0bl5 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b5c752 l0bl5 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b5c753 l0bl5 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b5c754 l0bl5 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b5c755 l0bl5 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b5c756 l0bl5 vdd x756 x756b CELLD r1=900e3 r0=10000e3
xl0b5c757 l0bl5 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b5c758 l0bl5 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b5c759 l0bl5 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b5c760 l0bl5 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b5c761 l0bl5 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b5c762 l0bl5 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b5c763 l0bl5 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b5c764 l0bl5 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b5c765 l0bl5 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b5c766 l0bl5 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b5c767 l0bl5 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b5c768 l0bl5 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b5c769 l0bl5 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b5c770 l0bl5 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b5c771 l0bl5 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b5c772 l0bl5 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b5c773 l0bl5 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b5c774 l0bl5 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b5c775 l0bl5 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b5c776 l0bl5 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b5c777 l0bl5 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b5c778 l0bl5 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b5c779 l0bl5 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b5c780 l0bl5 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b5c781 l0bl5 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b5c782 l0bl5 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b5c783 l0bl5 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b6c0 l0bl6 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b6c1 l0bl6 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b6c2 l0bl6 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b6c3 l0bl6 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b6c4 l0bl6 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b6c5 l0bl6 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b6c6 l0bl6 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b6c7 l0bl6 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b6c8 l0bl6 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b6c9 l0bl6 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b6c10 l0bl6 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b6c11 l0bl6 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b6c12 l0bl6 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b6c13 l0bl6 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b6c14 l0bl6 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b6c15 l0bl6 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b6c16 l0bl6 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b6c17 l0bl6 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b6c18 l0bl6 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b6c19 l0bl6 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b6c20 l0bl6 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b6c21 l0bl6 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b6c22 l0bl6 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b6c23 l0bl6 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b6c24 l0bl6 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b6c25 l0bl6 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b6c26 l0bl6 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b6c27 l0bl6 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b6c28 l0bl6 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b6c29 l0bl6 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b6c30 l0bl6 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b6c31 l0bl6 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b6c32 l0bl6 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b6c33 l0bl6 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b6c34 l0bl6 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b6c35 l0bl6 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b6c36 l0bl6 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b6c37 l0bl6 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b6c38 l0bl6 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b6c39 l0bl6 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b6c40 l0bl6 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b6c41 l0bl6 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b6c42 l0bl6 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b6c43 l0bl6 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b6c44 l0bl6 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b6c45 l0bl6 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b6c46 l0bl6 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b6c47 l0bl6 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b6c48 l0bl6 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b6c49 l0bl6 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b6c50 l0bl6 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b6c51 l0bl6 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b6c52 l0bl6 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b6c53 l0bl6 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b6c54 l0bl6 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b6c55 l0bl6 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b6c56 l0bl6 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b6c57 l0bl6 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b6c58 l0bl6 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b6c59 l0bl6 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b6c60 l0bl6 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b6c61 l0bl6 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b6c62 l0bl6 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b6c63 l0bl6 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b6c64 l0bl6 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b6c65 l0bl6 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b6c66 l0bl6 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b6c67 l0bl6 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b6c68 l0bl6 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b6c69 l0bl6 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b6c70 l0bl6 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b6c71 l0bl6 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b6c72 l0bl6 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b6c73 l0bl6 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b6c74 l0bl6 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b6c75 l0bl6 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b6c76 l0bl6 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b6c77 l0bl6 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b6c78 l0bl6 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b6c79 l0bl6 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b6c80 l0bl6 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b6c81 l0bl6 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b6c82 l0bl6 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b6c83 l0bl6 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b6c84 l0bl6 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b6c85 l0bl6 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b6c86 l0bl6 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b6c87 l0bl6 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b6c88 l0bl6 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b6c89 l0bl6 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b6c90 l0bl6 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b6c91 l0bl6 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b6c92 l0bl6 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b6c93 l0bl6 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b6c94 l0bl6 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b6c95 l0bl6 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b6c96 l0bl6 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b6c97 l0bl6 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b6c98 l0bl6 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b6c99 l0bl6 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b6c100 l0bl6 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b6c101 l0bl6 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b6c102 l0bl6 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b6c103 l0bl6 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b6c104 l0bl6 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b6c105 l0bl6 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b6c106 l0bl6 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b6c107 l0bl6 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b6c108 l0bl6 vdd x108 x108b CELLD r1=10000e3 r0=900e3
xl0b6c109 l0bl6 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b6c110 l0bl6 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b6c111 l0bl6 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b6c112 l0bl6 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b6c113 l0bl6 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b6c114 l0bl6 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b6c115 l0bl6 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b6c116 l0bl6 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b6c117 l0bl6 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b6c118 l0bl6 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b6c119 l0bl6 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b6c120 l0bl6 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b6c121 l0bl6 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b6c122 l0bl6 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b6c123 l0bl6 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b6c124 l0bl6 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b6c125 l0bl6 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b6c126 l0bl6 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b6c127 l0bl6 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b6c128 l0bl6 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b6c129 l0bl6 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b6c130 l0bl6 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b6c131 l0bl6 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b6c132 l0bl6 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b6c133 l0bl6 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b6c134 l0bl6 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b6c135 l0bl6 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b6c136 l0bl6 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b6c137 l0bl6 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b6c138 l0bl6 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b6c139 l0bl6 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b6c140 l0bl6 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b6c141 l0bl6 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b6c142 l0bl6 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b6c143 l0bl6 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b6c144 l0bl6 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b6c145 l0bl6 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b6c146 l0bl6 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b6c147 l0bl6 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b6c148 l0bl6 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b6c149 l0bl6 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b6c150 l0bl6 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b6c151 l0bl6 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b6c152 l0bl6 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b6c153 l0bl6 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b6c154 l0bl6 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b6c155 l0bl6 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b6c156 l0bl6 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b6c157 l0bl6 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b6c158 l0bl6 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b6c159 l0bl6 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b6c160 l0bl6 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b6c161 l0bl6 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b6c162 l0bl6 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b6c163 l0bl6 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b6c164 l0bl6 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b6c165 l0bl6 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b6c166 l0bl6 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b6c167 l0bl6 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b6c168 l0bl6 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b6c169 l0bl6 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b6c170 l0bl6 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b6c171 l0bl6 vdd x171 x171b CELLD r1=10000e3 r0=900e3
xl0b6c172 l0bl6 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b6c173 l0bl6 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b6c174 l0bl6 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b6c175 l0bl6 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b6c176 l0bl6 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b6c177 l0bl6 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b6c178 l0bl6 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b6c179 l0bl6 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b6c180 l0bl6 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b6c181 l0bl6 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b6c182 l0bl6 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b6c183 l0bl6 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b6c184 l0bl6 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b6c185 l0bl6 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b6c186 l0bl6 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b6c187 l0bl6 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b6c188 l0bl6 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b6c189 l0bl6 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b6c190 l0bl6 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b6c191 l0bl6 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b6c192 l0bl6 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b6c193 l0bl6 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b6c194 l0bl6 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b6c195 l0bl6 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b6c196 l0bl6 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b6c197 l0bl6 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b6c198 l0bl6 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b6c199 l0bl6 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b6c200 l0bl6 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b6c201 l0bl6 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b6c202 l0bl6 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b6c203 l0bl6 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b6c204 l0bl6 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b6c205 l0bl6 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b6c206 l0bl6 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b6c207 l0bl6 vdd x207 x207b CELLD r1=900e3 r0=10000e3
xl0b6c208 l0bl6 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b6c209 l0bl6 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b6c210 l0bl6 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b6c211 l0bl6 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b6c212 l0bl6 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b6c213 l0bl6 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b6c214 l0bl6 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b6c215 l0bl6 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b6c216 l0bl6 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b6c217 l0bl6 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b6c218 l0bl6 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b6c219 l0bl6 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b6c220 l0bl6 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b6c221 l0bl6 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b6c222 l0bl6 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b6c223 l0bl6 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b6c224 l0bl6 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b6c225 l0bl6 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b6c226 l0bl6 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b6c227 l0bl6 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b6c228 l0bl6 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b6c229 l0bl6 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b6c230 l0bl6 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b6c231 l0bl6 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b6c232 l0bl6 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b6c233 l0bl6 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b6c234 l0bl6 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b6c235 l0bl6 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b6c236 l0bl6 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b6c237 l0bl6 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b6c238 l0bl6 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b6c239 l0bl6 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b6c240 l0bl6 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b6c241 l0bl6 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b6c242 l0bl6 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b6c243 l0bl6 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b6c244 l0bl6 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b6c245 l0bl6 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b6c246 l0bl6 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b6c247 l0bl6 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b6c248 l0bl6 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b6c249 l0bl6 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b6c250 l0bl6 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b6c251 l0bl6 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b6c252 l0bl6 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b6c253 l0bl6 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b6c254 l0bl6 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b6c255 l0bl6 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b6c256 l0bl6 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b6c257 l0bl6 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b6c258 l0bl6 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b6c259 l0bl6 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b6c260 l0bl6 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b6c261 l0bl6 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b6c262 l0bl6 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b6c263 l0bl6 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b6c264 l0bl6 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b6c265 l0bl6 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b6c266 l0bl6 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b6c267 l0bl6 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b6c268 l0bl6 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b6c269 l0bl6 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b6c270 l0bl6 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b6c271 l0bl6 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b6c272 l0bl6 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b6c273 l0bl6 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b6c274 l0bl6 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b6c275 l0bl6 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b6c276 l0bl6 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b6c277 l0bl6 vdd x277 x277b CELLD r1=900e3 r0=10000e3
xl0b6c278 l0bl6 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b6c279 l0bl6 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b6c280 l0bl6 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b6c281 l0bl6 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b6c282 l0bl6 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b6c283 l0bl6 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b6c284 l0bl6 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b6c285 l0bl6 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b6c286 l0bl6 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b6c287 l0bl6 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b6c288 l0bl6 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b6c289 l0bl6 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b6c290 l0bl6 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b6c291 l0bl6 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b6c292 l0bl6 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b6c293 l0bl6 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b6c294 l0bl6 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b6c295 l0bl6 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b6c296 l0bl6 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b6c297 l0bl6 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b6c298 l0bl6 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b6c299 l0bl6 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b6c300 l0bl6 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b6c301 l0bl6 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b6c302 l0bl6 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b6c303 l0bl6 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b6c304 l0bl6 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b6c305 l0bl6 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b6c306 l0bl6 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b6c307 l0bl6 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b6c308 l0bl6 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b6c309 l0bl6 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b6c310 l0bl6 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b6c311 l0bl6 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b6c312 l0bl6 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b6c313 l0bl6 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b6c314 l0bl6 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b6c315 l0bl6 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b6c316 l0bl6 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b6c317 l0bl6 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b6c318 l0bl6 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b6c319 l0bl6 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b6c320 l0bl6 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b6c321 l0bl6 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b6c322 l0bl6 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b6c323 l0bl6 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b6c324 l0bl6 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b6c325 l0bl6 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b6c326 l0bl6 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b6c327 l0bl6 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b6c328 l0bl6 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b6c329 l0bl6 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b6c330 l0bl6 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b6c331 l0bl6 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b6c332 l0bl6 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b6c333 l0bl6 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b6c334 l0bl6 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b6c335 l0bl6 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b6c336 l0bl6 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b6c337 l0bl6 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b6c338 l0bl6 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b6c339 l0bl6 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b6c340 l0bl6 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b6c341 l0bl6 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b6c342 l0bl6 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b6c343 l0bl6 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b6c344 l0bl6 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b6c345 l0bl6 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b6c346 l0bl6 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b6c347 l0bl6 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b6c348 l0bl6 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b6c349 l0bl6 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b6c350 l0bl6 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b6c351 l0bl6 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b6c352 l0bl6 vdd x352 x352b CELLD r1=10000e3 r0=900e3
xl0b6c353 l0bl6 vdd x353 x353b CELLD r1=10000e3 r0=900e3
xl0b6c354 l0bl6 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b6c355 l0bl6 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b6c356 l0bl6 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b6c357 l0bl6 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b6c358 l0bl6 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b6c359 l0bl6 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b6c360 l0bl6 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b6c361 l0bl6 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b6c362 l0bl6 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b6c363 l0bl6 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b6c364 l0bl6 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b6c365 l0bl6 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b6c366 l0bl6 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b6c367 l0bl6 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b6c368 l0bl6 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b6c369 l0bl6 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b6c370 l0bl6 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b6c371 l0bl6 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b6c372 l0bl6 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b6c373 l0bl6 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b6c374 l0bl6 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b6c375 l0bl6 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b6c376 l0bl6 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b6c377 l0bl6 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b6c378 l0bl6 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b6c379 l0bl6 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b6c380 l0bl6 vdd x380 x380b CELLD r1=10000e3 r0=900e3
xl0b6c381 l0bl6 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b6c382 l0bl6 vdd x382 x382b CELLD r1=10000e3 r0=900e3
xl0b6c383 l0bl6 vdd x383 x383b CELLD r1=10000e3 r0=900e3
xl0b6c384 l0bl6 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b6c385 l0bl6 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b6c386 l0bl6 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b6c387 l0bl6 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b6c388 l0bl6 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b6c389 l0bl6 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b6c390 l0bl6 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b6c391 l0bl6 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b6c392 l0bl6 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b6c393 l0bl6 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b6c394 l0bl6 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b6c395 l0bl6 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b6c396 l0bl6 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b6c397 l0bl6 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b6c398 l0bl6 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b6c399 l0bl6 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b6c400 l0bl6 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b6c401 l0bl6 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b6c402 l0bl6 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b6c403 l0bl6 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b6c404 l0bl6 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b6c405 l0bl6 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b6c406 l0bl6 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b6c407 l0bl6 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b6c408 l0bl6 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b6c409 l0bl6 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b6c410 l0bl6 vdd x410 x410b CELLD r1=10000e3 r0=900e3
xl0b6c411 l0bl6 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b6c412 l0bl6 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b6c413 l0bl6 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b6c414 l0bl6 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b6c415 l0bl6 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b6c416 l0bl6 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b6c417 l0bl6 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b6c418 l0bl6 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b6c419 l0bl6 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b6c420 l0bl6 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b6c421 l0bl6 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b6c422 l0bl6 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b6c423 l0bl6 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b6c424 l0bl6 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b6c425 l0bl6 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b6c426 l0bl6 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b6c427 l0bl6 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b6c428 l0bl6 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b6c429 l0bl6 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b6c430 l0bl6 vdd x430 x430b CELLD r1=10000e3 r0=900e3
xl0b6c431 l0bl6 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b6c432 l0bl6 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b6c433 l0bl6 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b6c434 l0bl6 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b6c435 l0bl6 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b6c436 l0bl6 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b6c437 l0bl6 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b6c438 l0bl6 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b6c439 l0bl6 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b6c440 l0bl6 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b6c441 l0bl6 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b6c442 l0bl6 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b6c443 l0bl6 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b6c444 l0bl6 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b6c445 l0bl6 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b6c446 l0bl6 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b6c447 l0bl6 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b6c448 l0bl6 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b6c449 l0bl6 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b6c450 l0bl6 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b6c451 l0bl6 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b6c452 l0bl6 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b6c453 l0bl6 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b6c454 l0bl6 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b6c455 l0bl6 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b6c456 l0bl6 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b6c457 l0bl6 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b6c458 l0bl6 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b6c459 l0bl6 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b6c460 l0bl6 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b6c461 l0bl6 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b6c462 l0bl6 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b6c463 l0bl6 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b6c464 l0bl6 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b6c465 l0bl6 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b6c466 l0bl6 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b6c467 l0bl6 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b6c468 l0bl6 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b6c469 l0bl6 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b6c470 l0bl6 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b6c471 l0bl6 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b6c472 l0bl6 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b6c473 l0bl6 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b6c474 l0bl6 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b6c475 l0bl6 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b6c476 l0bl6 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b6c477 l0bl6 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b6c478 l0bl6 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b6c479 l0bl6 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b6c480 l0bl6 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b6c481 l0bl6 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b6c482 l0bl6 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b6c483 l0bl6 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b6c484 l0bl6 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b6c485 l0bl6 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b6c486 l0bl6 vdd x486 x486b CELLD r1=10000e3 r0=900e3
xl0b6c487 l0bl6 vdd x487 x487b CELLD r1=10000e3 r0=900e3
xl0b6c488 l0bl6 vdd x488 x488b CELLD r1=10000e3 r0=900e3
xl0b6c489 l0bl6 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b6c490 l0bl6 vdd x490 x490b CELLD r1=10000e3 r0=900e3
xl0b6c491 l0bl6 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b6c492 l0bl6 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b6c493 l0bl6 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b6c494 l0bl6 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b6c495 l0bl6 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b6c496 l0bl6 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b6c497 l0bl6 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b6c498 l0bl6 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b6c499 l0bl6 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b6c500 l0bl6 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b6c501 l0bl6 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b6c502 l0bl6 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b6c503 l0bl6 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b6c504 l0bl6 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b6c505 l0bl6 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b6c506 l0bl6 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b6c507 l0bl6 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b6c508 l0bl6 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b6c509 l0bl6 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b6c510 l0bl6 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b6c511 l0bl6 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b6c512 l0bl6 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b6c513 l0bl6 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b6c514 l0bl6 vdd x514 x514b CELLD r1=10000e3 r0=900e3
xl0b6c515 l0bl6 vdd x515 x515b CELLD r1=10000e3 r0=900e3
xl0b6c516 l0bl6 vdd x516 x516b CELLD r1=10000e3 r0=900e3
xl0b6c517 l0bl6 vdd x517 x517b CELLD r1=10000e3 r0=900e3
xl0b6c518 l0bl6 vdd x518 x518b CELLD r1=10000e3 r0=900e3
xl0b6c519 l0bl6 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b6c520 l0bl6 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b6c521 l0bl6 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b6c522 l0bl6 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b6c523 l0bl6 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b6c524 l0bl6 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b6c525 l0bl6 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b6c526 l0bl6 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b6c527 l0bl6 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b6c528 l0bl6 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b6c529 l0bl6 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b6c530 l0bl6 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b6c531 l0bl6 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b6c532 l0bl6 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b6c533 l0bl6 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b6c534 l0bl6 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b6c535 l0bl6 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b6c536 l0bl6 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b6c537 l0bl6 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b6c538 l0bl6 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b6c539 l0bl6 vdd x539 x539b CELLD r1=900e3 r0=10000e3
xl0b6c540 l0bl6 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b6c541 l0bl6 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b6c542 l0bl6 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b6c543 l0bl6 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b6c544 l0bl6 vdd x544 x544b CELLD r1=10000e3 r0=900e3
xl0b6c545 l0bl6 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b6c546 l0bl6 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b6c547 l0bl6 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b6c548 l0bl6 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b6c549 l0bl6 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b6c550 l0bl6 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b6c551 l0bl6 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b6c552 l0bl6 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b6c553 l0bl6 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b6c554 l0bl6 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b6c555 l0bl6 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b6c556 l0bl6 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b6c557 l0bl6 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b6c558 l0bl6 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b6c559 l0bl6 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b6c560 l0bl6 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b6c561 l0bl6 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b6c562 l0bl6 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b6c563 l0bl6 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b6c564 l0bl6 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b6c565 l0bl6 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b6c566 l0bl6 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b6c567 l0bl6 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b6c568 l0bl6 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b6c569 l0bl6 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b6c570 l0bl6 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b6c571 l0bl6 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b6c572 l0bl6 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b6c573 l0bl6 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b6c574 l0bl6 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b6c575 l0bl6 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b6c576 l0bl6 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b6c577 l0bl6 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b6c578 l0bl6 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b6c579 l0bl6 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b6c580 l0bl6 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b6c581 l0bl6 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b6c582 l0bl6 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b6c583 l0bl6 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b6c584 l0bl6 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b6c585 l0bl6 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b6c586 l0bl6 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b6c587 l0bl6 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b6c588 l0bl6 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b6c589 l0bl6 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b6c590 l0bl6 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b6c591 l0bl6 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b6c592 l0bl6 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b6c593 l0bl6 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b6c594 l0bl6 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b6c595 l0bl6 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b6c596 l0bl6 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b6c597 l0bl6 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b6c598 l0bl6 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b6c599 l0bl6 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b6c600 l0bl6 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b6c601 l0bl6 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b6c602 l0bl6 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b6c603 l0bl6 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b6c604 l0bl6 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b6c605 l0bl6 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b6c606 l0bl6 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b6c607 l0bl6 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b6c608 l0bl6 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b6c609 l0bl6 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b6c610 l0bl6 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b6c611 l0bl6 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b6c612 l0bl6 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b6c613 l0bl6 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b6c614 l0bl6 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b6c615 l0bl6 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b6c616 l0bl6 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b6c617 l0bl6 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b6c618 l0bl6 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b6c619 l0bl6 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b6c620 l0bl6 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b6c621 l0bl6 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b6c622 l0bl6 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b6c623 l0bl6 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b6c624 l0bl6 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b6c625 l0bl6 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b6c626 l0bl6 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b6c627 l0bl6 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b6c628 l0bl6 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b6c629 l0bl6 vdd x629 x629b CELLD r1=900e3 r0=10000e3
xl0b6c630 l0bl6 vdd x630 x630b CELLD r1=900e3 r0=10000e3
xl0b6c631 l0bl6 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b6c632 l0bl6 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b6c633 l0bl6 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b6c634 l0bl6 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b6c635 l0bl6 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b6c636 l0bl6 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b6c637 l0bl6 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b6c638 l0bl6 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b6c639 l0bl6 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b6c640 l0bl6 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b6c641 l0bl6 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b6c642 l0bl6 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b6c643 l0bl6 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b6c644 l0bl6 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b6c645 l0bl6 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b6c646 l0bl6 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b6c647 l0bl6 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b6c648 l0bl6 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b6c649 l0bl6 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b6c650 l0bl6 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b6c651 l0bl6 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b6c652 l0bl6 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b6c653 l0bl6 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b6c654 l0bl6 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b6c655 l0bl6 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b6c656 l0bl6 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b6c657 l0bl6 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b6c658 l0bl6 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b6c659 l0bl6 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b6c660 l0bl6 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b6c661 l0bl6 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b6c662 l0bl6 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b6c663 l0bl6 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b6c664 l0bl6 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b6c665 l0bl6 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b6c666 l0bl6 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b6c667 l0bl6 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b6c668 l0bl6 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b6c669 l0bl6 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b6c670 l0bl6 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b6c671 l0bl6 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b6c672 l0bl6 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b6c673 l0bl6 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b6c674 l0bl6 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b6c675 l0bl6 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b6c676 l0bl6 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b6c677 l0bl6 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b6c678 l0bl6 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b6c679 l0bl6 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b6c680 l0bl6 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b6c681 l0bl6 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b6c682 l0bl6 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b6c683 l0bl6 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b6c684 l0bl6 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b6c685 l0bl6 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b6c686 l0bl6 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b6c687 l0bl6 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b6c688 l0bl6 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b6c689 l0bl6 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b6c690 l0bl6 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b6c691 l0bl6 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b6c692 l0bl6 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b6c693 l0bl6 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b6c694 l0bl6 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b6c695 l0bl6 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b6c696 l0bl6 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b6c697 l0bl6 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b6c698 l0bl6 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b6c699 l0bl6 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b6c700 l0bl6 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b6c701 l0bl6 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b6c702 l0bl6 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b6c703 l0bl6 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b6c704 l0bl6 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b6c705 l0bl6 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b6c706 l0bl6 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b6c707 l0bl6 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b6c708 l0bl6 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b6c709 l0bl6 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b6c710 l0bl6 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b6c711 l0bl6 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b6c712 l0bl6 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b6c713 l0bl6 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b6c714 l0bl6 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b6c715 l0bl6 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b6c716 l0bl6 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b6c717 l0bl6 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b6c718 l0bl6 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b6c719 l0bl6 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b6c720 l0bl6 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b6c721 l0bl6 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b6c722 l0bl6 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b6c723 l0bl6 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b6c724 l0bl6 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b6c725 l0bl6 vdd x725 x725b CELLD r1=10000e3 r0=900e3
xl0b6c726 l0bl6 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b6c727 l0bl6 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b6c728 l0bl6 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b6c729 l0bl6 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b6c730 l0bl6 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b6c731 l0bl6 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b6c732 l0bl6 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b6c733 l0bl6 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b6c734 l0bl6 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b6c735 l0bl6 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b6c736 l0bl6 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b6c737 l0bl6 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b6c738 l0bl6 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b6c739 l0bl6 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b6c740 l0bl6 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b6c741 l0bl6 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b6c742 l0bl6 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b6c743 l0bl6 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b6c744 l0bl6 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b6c745 l0bl6 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b6c746 l0bl6 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b6c747 l0bl6 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b6c748 l0bl6 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b6c749 l0bl6 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b6c750 l0bl6 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b6c751 l0bl6 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b6c752 l0bl6 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b6c753 l0bl6 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b6c754 l0bl6 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b6c755 l0bl6 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b6c756 l0bl6 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b6c757 l0bl6 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b6c758 l0bl6 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b6c759 l0bl6 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b6c760 l0bl6 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b6c761 l0bl6 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b6c762 l0bl6 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b6c763 l0bl6 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b6c764 l0bl6 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b6c765 l0bl6 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b6c766 l0bl6 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b6c767 l0bl6 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b6c768 l0bl6 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b6c769 l0bl6 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b6c770 l0bl6 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b6c771 l0bl6 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b6c772 l0bl6 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b6c773 l0bl6 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b6c774 l0bl6 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b6c775 l0bl6 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b6c776 l0bl6 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b6c777 l0bl6 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b6c778 l0bl6 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b6c779 l0bl6 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b6c780 l0bl6 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b6c781 l0bl6 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b6c782 l0bl6 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b6c783 l0bl6 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b7c0 l0bl7 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b7c1 l0bl7 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b7c2 l0bl7 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b7c3 l0bl7 vdd x3 x3b CELLD r1=10000e3 r0=900e3
xl0b7c4 l0bl7 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b7c5 l0bl7 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b7c6 l0bl7 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b7c7 l0bl7 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b7c8 l0bl7 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b7c9 l0bl7 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b7c10 l0bl7 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b7c11 l0bl7 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b7c12 l0bl7 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b7c13 l0bl7 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b7c14 l0bl7 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b7c15 l0bl7 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b7c16 l0bl7 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b7c17 l0bl7 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b7c18 l0bl7 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b7c19 l0bl7 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b7c20 l0bl7 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b7c21 l0bl7 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b7c22 l0bl7 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b7c23 l0bl7 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b7c24 l0bl7 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b7c25 l0bl7 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b7c26 l0bl7 vdd x26 x26b CELLD r1=10000e3 r0=900e3
xl0b7c27 l0bl7 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b7c28 l0bl7 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b7c29 l0bl7 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b7c30 l0bl7 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b7c31 l0bl7 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b7c32 l0bl7 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b7c33 l0bl7 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b7c34 l0bl7 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b7c35 l0bl7 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b7c36 l0bl7 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b7c37 l0bl7 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b7c38 l0bl7 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b7c39 l0bl7 vdd x39 x39b CELLD r1=10000e3 r0=900e3
xl0b7c40 l0bl7 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b7c41 l0bl7 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b7c42 l0bl7 vdd x42 x42b CELLD r1=10000e3 r0=900e3
xl0b7c43 l0bl7 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b7c44 l0bl7 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b7c45 l0bl7 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b7c46 l0bl7 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b7c47 l0bl7 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b7c48 l0bl7 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b7c49 l0bl7 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b7c50 l0bl7 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b7c51 l0bl7 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b7c52 l0bl7 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b7c53 l0bl7 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b7c54 l0bl7 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b7c55 l0bl7 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b7c56 l0bl7 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b7c57 l0bl7 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b7c58 l0bl7 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b7c59 l0bl7 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b7c60 l0bl7 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b7c61 l0bl7 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b7c62 l0bl7 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b7c63 l0bl7 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b7c64 l0bl7 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b7c65 l0bl7 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b7c66 l0bl7 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b7c67 l0bl7 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b7c68 l0bl7 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b7c69 l0bl7 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b7c70 l0bl7 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b7c71 l0bl7 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b7c72 l0bl7 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b7c73 l0bl7 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b7c74 l0bl7 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b7c75 l0bl7 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b7c76 l0bl7 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b7c77 l0bl7 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b7c78 l0bl7 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b7c79 l0bl7 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b7c80 l0bl7 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b7c81 l0bl7 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b7c82 l0bl7 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b7c83 l0bl7 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b7c84 l0bl7 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b7c85 l0bl7 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b7c86 l0bl7 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b7c87 l0bl7 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b7c88 l0bl7 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b7c89 l0bl7 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b7c90 l0bl7 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b7c91 l0bl7 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b7c92 l0bl7 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b7c93 l0bl7 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b7c94 l0bl7 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b7c95 l0bl7 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b7c96 l0bl7 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b7c97 l0bl7 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b7c98 l0bl7 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b7c99 l0bl7 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b7c100 l0bl7 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b7c101 l0bl7 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b7c102 l0bl7 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b7c103 l0bl7 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b7c104 l0bl7 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b7c105 l0bl7 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b7c106 l0bl7 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b7c107 l0bl7 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b7c108 l0bl7 vdd x108 x108b CELLD r1=10000e3 r0=900e3
xl0b7c109 l0bl7 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b7c110 l0bl7 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b7c111 l0bl7 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b7c112 l0bl7 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b7c113 l0bl7 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b7c114 l0bl7 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b7c115 l0bl7 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b7c116 l0bl7 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b7c117 l0bl7 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b7c118 l0bl7 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b7c119 l0bl7 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b7c120 l0bl7 vdd x120 x120b CELLD r1=900e3 r0=10000e3
xl0b7c121 l0bl7 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b7c122 l0bl7 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b7c123 l0bl7 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b7c124 l0bl7 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b7c125 l0bl7 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b7c126 l0bl7 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b7c127 l0bl7 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b7c128 l0bl7 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b7c129 l0bl7 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b7c130 l0bl7 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b7c131 l0bl7 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b7c132 l0bl7 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b7c133 l0bl7 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b7c134 l0bl7 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b7c135 l0bl7 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b7c136 l0bl7 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b7c137 l0bl7 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b7c138 l0bl7 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b7c139 l0bl7 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b7c140 l0bl7 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b7c141 l0bl7 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b7c142 l0bl7 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b7c143 l0bl7 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b7c144 l0bl7 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b7c145 l0bl7 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b7c146 l0bl7 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b7c147 l0bl7 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b7c148 l0bl7 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b7c149 l0bl7 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b7c150 l0bl7 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b7c151 l0bl7 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b7c152 l0bl7 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b7c153 l0bl7 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b7c154 l0bl7 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b7c155 l0bl7 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b7c156 l0bl7 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b7c157 l0bl7 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b7c158 l0bl7 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b7c159 l0bl7 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b7c160 l0bl7 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b7c161 l0bl7 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b7c162 l0bl7 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b7c163 l0bl7 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b7c164 l0bl7 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b7c165 l0bl7 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b7c166 l0bl7 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b7c167 l0bl7 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b7c168 l0bl7 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b7c169 l0bl7 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b7c170 l0bl7 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b7c171 l0bl7 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b7c172 l0bl7 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b7c173 l0bl7 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b7c174 l0bl7 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b7c175 l0bl7 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b7c176 l0bl7 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b7c177 l0bl7 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b7c178 l0bl7 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b7c179 l0bl7 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b7c180 l0bl7 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b7c181 l0bl7 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b7c182 l0bl7 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b7c183 l0bl7 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b7c184 l0bl7 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b7c185 l0bl7 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b7c186 l0bl7 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b7c187 l0bl7 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b7c188 l0bl7 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b7c189 l0bl7 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b7c190 l0bl7 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b7c191 l0bl7 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b7c192 l0bl7 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b7c193 l0bl7 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b7c194 l0bl7 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b7c195 l0bl7 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b7c196 l0bl7 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b7c197 l0bl7 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b7c198 l0bl7 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b7c199 l0bl7 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b7c200 l0bl7 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b7c201 l0bl7 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b7c202 l0bl7 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b7c203 l0bl7 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b7c204 l0bl7 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b7c205 l0bl7 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b7c206 l0bl7 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b7c207 l0bl7 vdd x207 x207b CELLD r1=900e3 r0=10000e3
xl0b7c208 l0bl7 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b7c209 l0bl7 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b7c210 l0bl7 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b7c211 l0bl7 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b7c212 l0bl7 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b7c213 l0bl7 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b7c214 l0bl7 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b7c215 l0bl7 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b7c216 l0bl7 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b7c217 l0bl7 vdd x217 x217b CELLD r1=900e3 r0=10000e3
xl0b7c218 l0bl7 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b7c219 l0bl7 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b7c220 l0bl7 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b7c221 l0bl7 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b7c222 l0bl7 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b7c223 l0bl7 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b7c224 l0bl7 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b7c225 l0bl7 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b7c226 l0bl7 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b7c227 l0bl7 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b7c228 l0bl7 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b7c229 l0bl7 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b7c230 l0bl7 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b7c231 l0bl7 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b7c232 l0bl7 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b7c233 l0bl7 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b7c234 l0bl7 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b7c235 l0bl7 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b7c236 l0bl7 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b7c237 l0bl7 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b7c238 l0bl7 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b7c239 l0bl7 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b7c240 l0bl7 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b7c241 l0bl7 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b7c242 l0bl7 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b7c243 l0bl7 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b7c244 l0bl7 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b7c245 l0bl7 vdd x245 x245b CELLD r1=900e3 r0=10000e3
xl0b7c246 l0bl7 vdd x246 x246b CELLD r1=900e3 r0=10000e3
xl0b7c247 l0bl7 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b7c248 l0bl7 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b7c249 l0bl7 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b7c250 l0bl7 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b7c251 l0bl7 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b7c252 l0bl7 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b7c253 l0bl7 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b7c254 l0bl7 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b7c255 l0bl7 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b7c256 l0bl7 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b7c257 l0bl7 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b7c258 l0bl7 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b7c259 l0bl7 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b7c260 l0bl7 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b7c261 l0bl7 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b7c262 l0bl7 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b7c263 l0bl7 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b7c264 l0bl7 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b7c265 l0bl7 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b7c266 l0bl7 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b7c267 l0bl7 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b7c268 l0bl7 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b7c269 l0bl7 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b7c270 l0bl7 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b7c271 l0bl7 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b7c272 l0bl7 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b7c273 l0bl7 vdd x273 x273b CELLD r1=900e3 r0=10000e3
xl0b7c274 l0bl7 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b7c275 l0bl7 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b7c276 l0bl7 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b7c277 l0bl7 vdd x277 x277b CELLD r1=900e3 r0=10000e3
xl0b7c278 l0bl7 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b7c279 l0bl7 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b7c280 l0bl7 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b7c281 l0bl7 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b7c282 l0bl7 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b7c283 l0bl7 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b7c284 l0bl7 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b7c285 l0bl7 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b7c286 l0bl7 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b7c287 l0bl7 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b7c288 l0bl7 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b7c289 l0bl7 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b7c290 l0bl7 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b7c291 l0bl7 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b7c292 l0bl7 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b7c293 l0bl7 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b7c294 l0bl7 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b7c295 l0bl7 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b7c296 l0bl7 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b7c297 l0bl7 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b7c298 l0bl7 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b7c299 l0bl7 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b7c300 l0bl7 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b7c301 l0bl7 vdd x301 x301b CELLD r1=900e3 r0=10000e3
xl0b7c302 l0bl7 vdd x302 x302b CELLD r1=900e3 r0=10000e3
xl0b7c303 l0bl7 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b7c304 l0bl7 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b7c305 l0bl7 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b7c306 l0bl7 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b7c307 l0bl7 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b7c308 l0bl7 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b7c309 l0bl7 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b7c310 l0bl7 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b7c311 l0bl7 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b7c312 l0bl7 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b7c313 l0bl7 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b7c314 l0bl7 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b7c315 l0bl7 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b7c316 l0bl7 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b7c317 l0bl7 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b7c318 l0bl7 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b7c319 l0bl7 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b7c320 l0bl7 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b7c321 l0bl7 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b7c322 l0bl7 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b7c323 l0bl7 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b7c324 l0bl7 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b7c325 l0bl7 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b7c326 l0bl7 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b7c327 l0bl7 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b7c328 l0bl7 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b7c329 l0bl7 vdd x329 x329b CELLD r1=900e3 r0=10000e3
xl0b7c330 l0bl7 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b7c331 l0bl7 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b7c332 l0bl7 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b7c333 l0bl7 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b7c334 l0bl7 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b7c335 l0bl7 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b7c336 l0bl7 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b7c337 l0bl7 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b7c338 l0bl7 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b7c339 l0bl7 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b7c340 l0bl7 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b7c341 l0bl7 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b7c342 l0bl7 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b7c343 l0bl7 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b7c344 l0bl7 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b7c345 l0bl7 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b7c346 l0bl7 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b7c347 l0bl7 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b7c348 l0bl7 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b7c349 l0bl7 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b7c350 l0bl7 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b7c351 l0bl7 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b7c352 l0bl7 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b7c353 l0bl7 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b7c354 l0bl7 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b7c355 l0bl7 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b7c356 l0bl7 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b7c357 l0bl7 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b7c358 l0bl7 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b7c359 l0bl7 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b7c360 l0bl7 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b7c361 l0bl7 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b7c362 l0bl7 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b7c363 l0bl7 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b7c364 l0bl7 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b7c365 l0bl7 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b7c366 l0bl7 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b7c367 l0bl7 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b7c368 l0bl7 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b7c369 l0bl7 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b7c370 l0bl7 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b7c371 l0bl7 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b7c372 l0bl7 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b7c373 l0bl7 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b7c374 l0bl7 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b7c375 l0bl7 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b7c376 l0bl7 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b7c377 l0bl7 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b7c378 l0bl7 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b7c379 l0bl7 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b7c380 l0bl7 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b7c381 l0bl7 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b7c382 l0bl7 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b7c383 l0bl7 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b7c384 l0bl7 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b7c385 l0bl7 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b7c386 l0bl7 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b7c387 l0bl7 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b7c388 l0bl7 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b7c389 l0bl7 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b7c390 l0bl7 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b7c391 l0bl7 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b7c392 l0bl7 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b7c393 l0bl7 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b7c394 l0bl7 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b7c395 l0bl7 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b7c396 l0bl7 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b7c397 l0bl7 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b7c398 l0bl7 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b7c399 l0bl7 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b7c400 l0bl7 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b7c401 l0bl7 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b7c402 l0bl7 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b7c403 l0bl7 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b7c404 l0bl7 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b7c405 l0bl7 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b7c406 l0bl7 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b7c407 l0bl7 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b7c408 l0bl7 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b7c409 l0bl7 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b7c410 l0bl7 vdd x410 x410b CELLD r1=10000e3 r0=900e3
xl0b7c411 l0bl7 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b7c412 l0bl7 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b7c413 l0bl7 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b7c414 l0bl7 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b7c415 l0bl7 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b7c416 l0bl7 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b7c417 l0bl7 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b7c418 l0bl7 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b7c419 l0bl7 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b7c420 l0bl7 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b7c421 l0bl7 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b7c422 l0bl7 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b7c423 l0bl7 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b7c424 l0bl7 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b7c425 l0bl7 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b7c426 l0bl7 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b7c427 l0bl7 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b7c428 l0bl7 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b7c429 l0bl7 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b7c430 l0bl7 vdd x430 x430b CELLD r1=10000e3 r0=900e3
xl0b7c431 l0bl7 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b7c432 l0bl7 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b7c433 l0bl7 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b7c434 l0bl7 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b7c435 l0bl7 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b7c436 l0bl7 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b7c437 l0bl7 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b7c438 l0bl7 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b7c439 l0bl7 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b7c440 l0bl7 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b7c441 l0bl7 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b7c442 l0bl7 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b7c443 l0bl7 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b7c444 l0bl7 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b7c445 l0bl7 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b7c446 l0bl7 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b7c447 l0bl7 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b7c448 l0bl7 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b7c449 l0bl7 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b7c450 l0bl7 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b7c451 l0bl7 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b7c452 l0bl7 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b7c453 l0bl7 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b7c454 l0bl7 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b7c455 l0bl7 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b7c456 l0bl7 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b7c457 l0bl7 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b7c458 l0bl7 vdd x458 x458b CELLD r1=10000e3 r0=900e3
xl0b7c459 l0bl7 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b7c460 l0bl7 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b7c461 l0bl7 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b7c462 l0bl7 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b7c463 l0bl7 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b7c464 l0bl7 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b7c465 l0bl7 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b7c466 l0bl7 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b7c467 l0bl7 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b7c468 l0bl7 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b7c469 l0bl7 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b7c470 l0bl7 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b7c471 l0bl7 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b7c472 l0bl7 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b7c473 l0bl7 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b7c474 l0bl7 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b7c475 l0bl7 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b7c476 l0bl7 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b7c477 l0bl7 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b7c478 l0bl7 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b7c479 l0bl7 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b7c480 l0bl7 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b7c481 l0bl7 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b7c482 l0bl7 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b7c483 l0bl7 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b7c484 l0bl7 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b7c485 l0bl7 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b7c486 l0bl7 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b7c487 l0bl7 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b7c488 l0bl7 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b7c489 l0bl7 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b7c490 l0bl7 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b7c491 l0bl7 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b7c492 l0bl7 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b7c493 l0bl7 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b7c494 l0bl7 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b7c495 l0bl7 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b7c496 l0bl7 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b7c497 l0bl7 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b7c498 l0bl7 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b7c499 l0bl7 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b7c500 l0bl7 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b7c501 l0bl7 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b7c502 l0bl7 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b7c503 l0bl7 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b7c504 l0bl7 vdd x504 x504b CELLD r1=10000e3 r0=900e3
xl0b7c505 l0bl7 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b7c506 l0bl7 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b7c507 l0bl7 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b7c508 l0bl7 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b7c509 l0bl7 vdd x509 x509b CELLD r1=900e3 r0=10000e3
xl0b7c510 l0bl7 vdd x510 x510b CELLD r1=900e3 r0=10000e3
xl0b7c511 l0bl7 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b7c512 l0bl7 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b7c513 l0bl7 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b7c514 l0bl7 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b7c515 l0bl7 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b7c516 l0bl7 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b7c517 l0bl7 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b7c518 l0bl7 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b7c519 l0bl7 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b7c520 l0bl7 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b7c521 l0bl7 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b7c522 l0bl7 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b7c523 l0bl7 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b7c524 l0bl7 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b7c525 l0bl7 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b7c526 l0bl7 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b7c527 l0bl7 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b7c528 l0bl7 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b7c529 l0bl7 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b7c530 l0bl7 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b7c531 l0bl7 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b7c532 l0bl7 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b7c533 l0bl7 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b7c534 l0bl7 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b7c535 l0bl7 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b7c536 l0bl7 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b7c537 l0bl7 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b7c538 l0bl7 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b7c539 l0bl7 vdd x539 x539b CELLD r1=900e3 r0=10000e3
xl0b7c540 l0bl7 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b7c541 l0bl7 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b7c542 l0bl7 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b7c543 l0bl7 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b7c544 l0bl7 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b7c545 l0bl7 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b7c546 l0bl7 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b7c547 l0bl7 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b7c548 l0bl7 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b7c549 l0bl7 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b7c550 l0bl7 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b7c551 l0bl7 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b7c552 l0bl7 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b7c553 l0bl7 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b7c554 l0bl7 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b7c555 l0bl7 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b7c556 l0bl7 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b7c557 l0bl7 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b7c558 l0bl7 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b7c559 l0bl7 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b7c560 l0bl7 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b7c561 l0bl7 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b7c562 l0bl7 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b7c563 l0bl7 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b7c564 l0bl7 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b7c565 l0bl7 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b7c566 l0bl7 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b7c567 l0bl7 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b7c568 l0bl7 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b7c569 l0bl7 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b7c570 l0bl7 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b7c571 l0bl7 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b7c572 l0bl7 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b7c573 l0bl7 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b7c574 l0bl7 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b7c575 l0bl7 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b7c576 l0bl7 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b7c577 l0bl7 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b7c578 l0bl7 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b7c579 l0bl7 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b7c580 l0bl7 vdd x580 x580b CELLD r1=900e3 r0=10000e3
xl0b7c581 l0bl7 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b7c582 l0bl7 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b7c583 l0bl7 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b7c584 l0bl7 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b7c585 l0bl7 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b7c586 l0bl7 vdd x586 x586b CELLD r1=10000e3 r0=900e3
xl0b7c587 l0bl7 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b7c588 l0bl7 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b7c589 l0bl7 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b7c590 l0bl7 vdd x590 x590b CELLD r1=10000e3 r0=900e3
xl0b7c591 l0bl7 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b7c592 l0bl7 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b7c593 l0bl7 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b7c594 l0bl7 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b7c595 l0bl7 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b7c596 l0bl7 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b7c597 l0bl7 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b7c598 l0bl7 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b7c599 l0bl7 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b7c600 l0bl7 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b7c601 l0bl7 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b7c602 l0bl7 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b7c603 l0bl7 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b7c604 l0bl7 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b7c605 l0bl7 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b7c606 l0bl7 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b7c607 l0bl7 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b7c608 l0bl7 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b7c609 l0bl7 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b7c610 l0bl7 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b7c611 l0bl7 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b7c612 l0bl7 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b7c613 l0bl7 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b7c614 l0bl7 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b7c615 l0bl7 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b7c616 l0bl7 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b7c617 l0bl7 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b7c618 l0bl7 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b7c619 l0bl7 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b7c620 l0bl7 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b7c621 l0bl7 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b7c622 l0bl7 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b7c623 l0bl7 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b7c624 l0bl7 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b7c625 l0bl7 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b7c626 l0bl7 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b7c627 l0bl7 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b7c628 l0bl7 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b7c629 l0bl7 vdd x629 x629b CELLD r1=900e3 r0=10000e3
xl0b7c630 l0bl7 vdd x630 x630b CELLD r1=900e3 r0=10000e3
xl0b7c631 l0bl7 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b7c632 l0bl7 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b7c633 l0bl7 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b7c634 l0bl7 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b7c635 l0bl7 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b7c636 l0bl7 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b7c637 l0bl7 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b7c638 l0bl7 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b7c639 l0bl7 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b7c640 l0bl7 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b7c641 l0bl7 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b7c642 l0bl7 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b7c643 l0bl7 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b7c644 l0bl7 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b7c645 l0bl7 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b7c646 l0bl7 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b7c647 l0bl7 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b7c648 l0bl7 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b7c649 l0bl7 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b7c650 l0bl7 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b7c651 l0bl7 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b7c652 l0bl7 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b7c653 l0bl7 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b7c654 l0bl7 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b7c655 l0bl7 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b7c656 l0bl7 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b7c657 l0bl7 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b7c658 l0bl7 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b7c659 l0bl7 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b7c660 l0bl7 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b7c661 l0bl7 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b7c662 l0bl7 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b7c663 l0bl7 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b7c664 l0bl7 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b7c665 l0bl7 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b7c666 l0bl7 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b7c667 l0bl7 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b7c668 l0bl7 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b7c669 l0bl7 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b7c670 l0bl7 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b7c671 l0bl7 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b7c672 l0bl7 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b7c673 l0bl7 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b7c674 l0bl7 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b7c675 l0bl7 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b7c676 l0bl7 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b7c677 l0bl7 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b7c678 l0bl7 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b7c679 l0bl7 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b7c680 l0bl7 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b7c681 l0bl7 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b7c682 l0bl7 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b7c683 l0bl7 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b7c684 l0bl7 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b7c685 l0bl7 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b7c686 l0bl7 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b7c687 l0bl7 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b7c688 l0bl7 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b7c689 l0bl7 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b7c690 l0bl7 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b7c691 l0bl7 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b7c692 l0bl7 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b7c693 l0bl7 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b7c694 l0bl7 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b7c695 l0bl7 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b7c696 l0bl7 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b7c697 l0bl7 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b7c698 l0bl7 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b7c699 l0bl7 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b7c700 l0bl7 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b7c701 l0bl7 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b7c702 l0bl7 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b7c703 l0bl7 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b7c704 l0bl7 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b7c705 l0bl7 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b7c706 l0bl7 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b7c707 l0bl7 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b7c708 l0bl7 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b7c709 l0bl7 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b7c710 l0bl7 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b7c711 l0bl7 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b7c712 l0bl7 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b7c713 l0bl7 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b7c714 l0bl7 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b7c715 l0bl7 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b7c716 l0bl7 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b7c717 l0bl7 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b7c718 l0bl7 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b7c719 l0bl7 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b7c720 l0bl7 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b7c721 l0bl7 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b7c722 l0bl7 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b7c723 l0bl7 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b7c724 l0bl7 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b7c725 l0bl7 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b7c726 l0bl7 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b7c727 l0bl7 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b7c728 l0bl7 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b7c729 l0bl7 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b7c730 l0bl7 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b7c731 l0bl7 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b7c732 l0bl7 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b7c733 l0bl7 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b7c734 l0bl7 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b7c735 l0bl7 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b7c736 l0bl7 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b7c737 l0bl7 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b7c738 l0bl7 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b7c739 l0bl7 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b7c740 l0bl7 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b7c741 l0bl7 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b7c742 l0bl7 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b7c743 l0bl7 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b7c744 l0bl7 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b7c745 l0bl7 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b7c746 l0bl7 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b7c747 l0bl7 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b7c748 l0bl7 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b7c749 l0bl7 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b7c750 l0bl7 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b7c751 l0bl7 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b7c752 l0bl7 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b7c753 l0bl7 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b7c754 l0bl7 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b7c755 l0bl7 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b7c756 l0bl7 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b7c757 l0bl7 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b7c758 l0bl7 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b7c759 l0bl7 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b7c760 l0bl7 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b7c761 l0bl7 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b7c762 l0bl7 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b7c763 l0bl7 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b7c764 l0bl7 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b7c765 l0bl7 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b7c766 l0bl7 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b7c767 l0bl7 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b7c768 l0bl7 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b7c769 l0bl7 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b7c770 l0bl7 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b7c771 l0bl7 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b7c772 l0bl7 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b7c773 l0bl7 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b7c774 l0bl7 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b7c775 l0bl7 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b7c776 l0bl7 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b7c777 l0bl7 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b7c778 l0bl7 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b7c779 l0bl7 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b7c780 l0bl7 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b7c781 l0bl7 vdd x781 x781b CELLD r1=10000e3 r0=900e3
xl0b7c782 l0bl7 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b7c783 l0bl7 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b8c0 l0bl8 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b8c1 l0bl8 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b8c2 l0bl8 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b8c3 l0bl8 vdd x3 x3b CELLD r1=10000e3 r0=900e3
xl0b8c4 l0bl8 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b8c5 l0bl8 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b8c6 l0bl8 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b8c7 l0bl8 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b8c8 l0bl8 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b8c9 l0bl8 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b8c10 l0bl8 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b8c11 l0bl8 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b8c12 l0bl8 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b8c13 l0bl8 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b8c14 l0bl8 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b8c15 l0bl8 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b8c16 l0bl8 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b8c17 l0bl8 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b8c18 l0bl8 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b8c19 l0bl8 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b8c20 l0bl8 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b8c21 l0bl8 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b8c22 l0bl8 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b8c23 l0bl8 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b8c24 l0bl8 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b8c25 l0bl8 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b8c26 l0bl8 vdd x26 x26b CELLD r1=10000e3 r0=900e3
xl0b8c27 l0bl8 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b8c28 l0bl8 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b8c29 l0bl8 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b8c30 l0bl8 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b8c31 l0bl8 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b8c32 l0bl8 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b8c33 l0bl8 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b8c34 l0bl8 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b8c35 l0bl8 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b8c36 l0bl8 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b8c37 l0bl8 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b8c38 l0bl8 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b8c39 l0bl8 vdd x39 x39b CELLD r1=10000e3 r0=900e3
xl0b8c40 l0bl8 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b8c41 l0bl8 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b8c42 l0bl8 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b8c43 l0bl8 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b8c44 l0bl8 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b8c45 l0bl8 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b8c46 l0bl8 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b8c47 l0bl8 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b8c48 l0bl8 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b8c49 l0bl8 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b8c50 l0bl8 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b8c51 l0bl8 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b8c52 l0bl8 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b8c53 l0bl8 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b8c54 l0bl8 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b8c55 l0bl8 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b8c56 l0bl8 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b8c57 l0bl8 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b8c58 l0bl8 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b8c59 l0bl8 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b8c60 l0bl8 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b8c61 l0bl8 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b8c62 l0bl8 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b8c63 l0bl8 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b8c64 l0bl8 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b8c65 l0bl8 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b8c66 l0bl8 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b8c67 l0bl8 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b8c68 l0bl8 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b8c69 l0bl8 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b8c70 l0bl8 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b8c71 l0bl8 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b8c72 l0bl8 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b8c73 l0bl8 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b8c74 l0bl8 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b8c75 l0bl8 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b8c76 l0bl8 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b8c77 l0bl8 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b8c78 l0bl8 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b8c79 l0bl8 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b8c80 l0bl8 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b8c81 l0bl8 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b8c82 l0bl8 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b8c83 l0bl8 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b8c84 l0bl8 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b8c85 l0bl8 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b8c86 l0bl8 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b8c87 l0bl8 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b8c88 l0bl8 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b8c89 l0bl8 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b8c90 l0bl8 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b8c91 l0bl8 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b8c92 l0bl8 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b8c93 l0bl8 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b8c94 l0bl8 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b8c95 l0bl8 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b8c96 l0bl8 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b8c97 l0bl8 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b8c98 l0bl8 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b8c99 l0bl8 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b8c100 l0bl8 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b8c101 l0bl8 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b8c102 l0bl8 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b8c103 l0bl8 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b8c104 l0bl8 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b8c105 l0bl8 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b8c106 l0bl8 vdd x106 x106b CELLD r1=10000e3 r0=900e3
xl0b8c107 l0bl8 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b8c108 l0bl8 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b8c109 l0bl8 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b8c110 l0bl8 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b8c111 l0bl8 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b8c112 l0bl8 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b8c113 l0bl8 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b8c114 l0bl8 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b8c115 l0bl8 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b8c116 l0bl8 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b8c117 l0bl8 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b8c118 l0bl8 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b8c119 l0bl8 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b8c120 l0bl8 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b8c121 l0bl8 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b8c122 l0bl8 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b8c123 l0bl8 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b8c124 l0bl8 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b8c125 l0bl8 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b8c126 l0bl8 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b8c127 l0bl8 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b8c128 l0bl8 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b8c129 l0bl8 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b8c130 l0bl8 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b8c131 l0bl8 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b8c132 l0bl8 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b8c133 l0bl8 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b8c134 l0bl8 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b8c135 l0bl8 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b8c136 l0bl8 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b8c137 l0bl8 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b8c138 l0bl8 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b8c139 l0bl8 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b8c140 l0bl8 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b8c141 l0bl8 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b8c142 l0bl8 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b8c143 l0bl8 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b8c144 l0bl8 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b8c145 l0bl8 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b8c146 l0bl8 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b8c147 l0bl8 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b8c148 l0bl8 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b8c149 l0bl8 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b8c150 l0bl8 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b8c151 l0bl8 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b8c152 l0bl8 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b8c153 l0bl8 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b8c154 l0bl8 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b8c155 l0bl8 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b8c156 l0bl8 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b8c157 l0bl8 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b8c158 l0bl8 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b8c159 l0bl8 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b8c160 l0bl8 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b8c161 l0bl8 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b8c162 l0bl8 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b8c163 l0bl8 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b8c164 l0bl8 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b8c165 l0bl8 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b8c166 l0bl8 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b8c167 l0bl8 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b8c168 l0bl8 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b8c169 l0bl8 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b8c170 l0bl8 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b8c171 l0bl8 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b8c172 l0bl8 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b8c173 l0bl8 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b8c174 l0bl8 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b8c175 l0bl8 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b8c176 l0bl8 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b8c177 l0bl8 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b8c178 l0bl8 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b8c179 l0bl8 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b8c180 l0bl8 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b8c181 l0bl8 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b8c182 l0bl8 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b8c183 l0bl8 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b8c184 l0bl8 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b8c185 l0bl8 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b8c186 l0bl8 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b8c187 l0bl8 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b8c188 l0bl8 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b8c189 l0bl8 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b8c190 l0bl8 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b8c191 l0bl8 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b8c192 l0bl8 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b8c193 l0bl8 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b8c194 l0bl8 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b8c195 l0bl8 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b8c196 l0bl8 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b8c197 l0bl8 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b8c198 l0bl8 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b8c199 l0bl8 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b8c200 l0bl8 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b8c201 l0bl8 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b8c202 l0bl8 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b8c203 l0bl8 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b8c204 l0bl8 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b8c205 l0bl8 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b8c206 l0bl8 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b8c207 l0bl8 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b8c208 l0bl8 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b8c209 l0bl8 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b8c210 l0bl8 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b8c211 l0bl8 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b8c212 l0bl8 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b8c213 l0bl8 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b8c214 l0bl8 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b8c215 l0bl8 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b8c216 l0bl8 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b8c217 l0bl8 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b8c218 l0bl8 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b8c219 l0bl8 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b8c220 l0bl8 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b8c221 l0bl8 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b8c222 l0bl8 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b8c223 l0bl8 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b8c224 l0bl8 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b8c225 l0bl8 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b8c226 l0bl8 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b8c227 l0bl8 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b8c228 l0bl8 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b8c229 l0bl8 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b8c230 l0bl8 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b8c231 l0bl8 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b8c232 l0bl8 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b8c233 l0bl8 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b8c234 l0bl8 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b8c235 l0bl8 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b8c236 l0bl8 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b8c237 l0bl8 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b8c238 l0bl8 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b8c239 l0bl8 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b8c240 l0bl8 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b8c241 l0bl8 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b8c242 l0bl8 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b8c243 l0bl8 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b8c244 l0bl8 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b8c245 l0bl8 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b8c246 l0bl8 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b8c247 l0bl8 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b8c248 l0bl8 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b8c249 l0bl8 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b8c250 l0bl8 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b8c251 l0bl8 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b8c252 l0bl8 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b8c253 l0bl8 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b8c254 l0bl8 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b8c255 l0bl8 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b8c256 l0bl8 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b8c257 l0bl8 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b8c258 l0bl8 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b8c259 l0bl8 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b8c260 l0bl8 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b8c261 l0bl8 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b8c262 l0bl8 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b8c263 l0bl8 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b8c264 l0bl8 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b8c265 l0bl8 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b8c266 l0bl8 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b8c267 l0bl8 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b8c268 l0bl8 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b8c269 l0bl8 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b8c270 l0bl8 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b8c271 l0bl8 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b8c272 l0bl8 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b8c273 l0bl8 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b8c274 l0bl8 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b8c275 l0bl8 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b8c276 l0bl8 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b8c277 l0bl8 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b8c278 l0bl8 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b8c279 l0bl8 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b8c280 l0bl8 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b8c281 l0bl8 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b8c282 l0bl8 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b8c283 l0bl8 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b8c284 l0bl8 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b8c285 l0bl8 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b8c286 l0bl8 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b8c287 l0bl8 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b8c288 l0bl8 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b8c289 l0bl8 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b8c290 l0bl8 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b8c291 l0bl8 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b8c292 l0bl8 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b8c293 l0bl8 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b8c294 l0bl8 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b8c295 l0bl8 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b8c296 l0bl8 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b8c297 l0bl8 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b8c298 l0bl8 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b8c299 l0bl8 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b8c300 l0bl8 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b8c301 l0bl8 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b8c302 l0bl8 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b8c303 l0bl8 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b8c304 l0bl8 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b8c305 l0bl8 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b8c306 l0bl8 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b8c307 l0bl8 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b8c308 l0bl8 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b8c309 l0bl8 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b8c310 l0bl8 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b8c311 l0bl8 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b8c312 l0bl8 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b8c313 l0bl8 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b8c314 l0bl8 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b8c315 l0bl8 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b8c316 l0bl8 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b8c317 l0bl8 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b8c318 l0bl8 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b8c319 l0bl8 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b8c320 l0bl8 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b8c321 l0bl8 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b8c322 l0bl8 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b8c323 l0bl8 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b8c324 l0bl8 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b8c325 l0bl8 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b8c326 l0bl8 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b8c327 l0bl8 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b8c328 l0bl8 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b8c329 l0bl8 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b8c330 l0bl8 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b8c331 l0bl8 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b8c332 l0bl8 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b8c333 l0bl8 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b8c334 l0bl8 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b8c335 l0bl8 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b8c336 l0bl8 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b8c337 l0bl8 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b8c338 l0bl8 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b8c339 l0bl8 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b8c340 l0bl8 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b8c341 l0bl8 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b8c342 l0bl8 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b8c343 l0bl8 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b8c344 l0bl8 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b8c345 l0bl8 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b8c346 l0bl8 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b8c347 l0bl8 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b8c348 l0bl8 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b8c349 l0bl8 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b8c350 l0bl8 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b8c351 l0bl8 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b8c352 l0bl8 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b8c353 l0bl8 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b8c354 l0bl8 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b8c355 l0bl8 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b8c356 l0bl8 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b8c357 l0bl8 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b8c358 l0bl8 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b8c359 l0bl8 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b8c360 l0bl8 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b8c361 l0bl8 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b8c362 l0bl8 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b8c363 l0bl8 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b8c364 l0bl8 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b8c365 l0bl8 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b8c366 l0bl8 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b8c367 l0bl8 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b8c368 l0bl8 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b8c369 l0bl8 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b8c370 l0bl8 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b8c371 l0bl8 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b8c372 l0bl8 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b8c373 l0bl8 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b8c374 l0bl8 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b8c375 l0bl8 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b8c376 l0bl8 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b8c377 l0bl8 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b8c378 l0bl8 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b8c379 l0bl8 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b8c380 l0bl8 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b8c381 l0bl8 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b8c382 l0bl8 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b8c383 l0bl8 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b8c384 l0bl8 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b8c385 l0bl8 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b8c386 l0bl8 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b8c387 l0bl8 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b8c388 l0bl8 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b8c389 l0bl8 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b8c390 l0bl8 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b8c391 l0bl8 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b8c392 l0bl8 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b8c393 l0bl8 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b8c394 l0bl8 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b8c395 l0bl8 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b8c396 l0bl8 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b8c397 l0bl8 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b8c398 l0bl8 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b8c399 l0bl8 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b8c400 l0bl8 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b8c401 l0bl8 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b8c402 l0bl8 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b8c403 l0bl8 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b8c404 l0bl8 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b8c405 l0bl8 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b8c406 l0bl8 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b8c407 l0bl8 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b8c408 l0bl8 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b8c409 l0bl8 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b8c410 l0bl8 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b8c411 l0bl8 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b8c412 l0bl8 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b8c413 l0bl8 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b8c414 l0bl8 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b8c415 l0bl8 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b8c416 l0bl8 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b8c417 l0bl8 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b8c418 l0bl8 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b8c419 l0bl8 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b8c420 l0bl8 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b8c421 l0bl8 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b8c422 l0bl8 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b8c423 l0bl8 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b8c424 l0bl8 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b8c425 l0bl8 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b8c426 l0bl8 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b8c427 l0bl8 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b8c428 l0bl8 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b8c429 l0bl8 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b8c430 l0bl8 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b8c431 l0bl8 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b8c432 l0bl8 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b8c433 l0bl8 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b8c434 l0bl8 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b8c435 l0bl8 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b8c436 l0bl8 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b8c437 l0bl8 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b8c438 l0bl8 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b8c439 l0bl8 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b8c440 l0bl8 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b8c441 l0bl8 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b8c442 l0bl8 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b8c443 l0bl8 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b8c444 l0bl8 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b8c445 l0bl8 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b8c446 l0bl8 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b8c447 l0bl8 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b8c448 l0bl8 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b8c449 l0bl8 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b8c450 l0bl8 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b8c451 l0bl8 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b8c452 l0bl8 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b8c453 l0bl8 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b8c454 l0bl8 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b8c455 l0bl8 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b8c456 l0bl8 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b8c457 l0bl8 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b8c458 l0bl8 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b8c459 l0bl8 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b8c460 l0bl8 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b8c461 l0bl8 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b8c462 l0bl8 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b8c463 l0bl8 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b8c464 l0bl8 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b8c465 l0bl8 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b8c466 l0bl8 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b8c467 l0bl8 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b8c468 l0bl8 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b8c469 l0bl8 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b8c470 l0bl8 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b8c471 l0bl8 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b8c472 l0bl8 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b8c473 l0bl8 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b8c474 l0bl8 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b8c475 l0bl8 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b8c476 l0bl8 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b8c477 l0bl8 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b8c478 l0bl8 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b8c479 l0bl8 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b8c480 l0bl8 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b8c481 l0bl8 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b8c482 l0bl8 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b8c483 l0bl8 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b8c484 l0bl8 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b8c485 l0bl8 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b8c486 l0bl8 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b8c487 l0bl8 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b8c488 l0bl8 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b8c489 l0bl8 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b8c490 l0bl8 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b8c491 l0bl8 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b8c492 l0bl8 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b8c493 l0bl8 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b8c494 l0bl8 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b8c495 l0bl8 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b8c496 l0bl8 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b8c497 l0bl8 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b8c498 l0bl8 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b8c499 l0bl8 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b8c500 l0bl8 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b8c501 l0bl8 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b8c502 l0bl8 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b8c503 l0bl8 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b8c504 l0bl8 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b8c505 l0bl8 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b8c506 l0bl8 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b8c507 l0bl8 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b8c508 l0bl8 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b8c509 l0bl8 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b8c510 l0bl8 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b8c511 l0bl8 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b8c512 l0bl8 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b8c513 l0bl8 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b8c514 l0bl8 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b8c515 l0bl8 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b8c516 l0bl8 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b8c517 l0bl8 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b8c518 l0bl8 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b8c519 l0bl8 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b8c520 l0bl8 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b8c521 l0bl8 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b8c522 l0bl8 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b8c523 l0bl8 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b8c524 l0bl8 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b8c525 l0bl8 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b8c526 l0bl8 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b8c527 l0bl8 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b8c528 l0bl8 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b8c529 l0bl8 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b8c530 l0bl8 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b8c531 l0bl8 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b8c532 l0bl8 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b8c533 l0bl8 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b8c534 l0bl8 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b8c535 l0bl8 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b8c536 l0bl8 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b8c537 l0bl8 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b8c538 l0bl8 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b8c539 l0bl8 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b8c540 l0bl8 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b8c541 l0bl8 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b8c542 l0bl8 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b8c543 l0bl8 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b8c544 l0bl8 vdd x544 x544b CELLD r1=10000e3 r0=900e3
xl0b8c545 l0bl8 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b8c546 l0bl8 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b8c547 l0bl8 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b8c548 l0bl8 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b8c549 l0bl8 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b8c550 l0bl8 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b8c551 l0bl8 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b8c552 l0bl8 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b8c553 l0bl8 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b8c554 l0bl8 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b8c555 l0bl8 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b8c556 l0bl8 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b8c557 l0bl8 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b8c558 l0bl8 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b8c559 l0bl8 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b8c560 l0bl8 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b8c561 l0bl8 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b8c562 l0bl8 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b8c563 l0bl8 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b8c564 l0bl8 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b8c565 l0bl8 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b8c566 l0bl8 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b8c567 l0bl8 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b8c568 l0bl8 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b8c569 l0bl8 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b8c570 l0bl8 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b8c571 l0bl8 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b8c572 l0bl8 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b8c573 l0bl8 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b8c574 l0bl8 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b8c575 l0bl8 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b8c576 l0bl8 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b8c577 l0bl8 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b8c578 l0bl8 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b8c579 l0bl8 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b8c580 l0bl8 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b8c581 l0bl8 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b8c582 l0bl8 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b8c583 l0bl8 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b8c584 l0bl8 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b8c585 l0bl8 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b8c586 l0bl8 vdd x586 x586b CELLD r1=10000e3 r0=900e3
xl0b8c587 l0bl8 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b8c588 l0bl8 vdd x588 x588b CELLD r1=10000e3 r0=900e3
xl0b8c589 l0bl8 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b8c590 l0bl8 vdd x590 x590b CELLD r1=10000e3 r0=900e3
xl0b8c591 l0bl8 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b8c592 l0bl8 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b8c593 l0bl8 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b8c594 l0bl8 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b8c595 l0bl8 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b8c596 l0bl8 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b8c597 l0bl8 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b8c598 l0bl8 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b8c599 l0bl8 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b8c600 l0bl8 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b8c601 l0bl8 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b8c602 l0bl8 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b8c603 l0bl8 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b8c604 l0bl8 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b8c605 l0bl8 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b8c606 l0bl8 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b8c607 l0bl8 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b8c608 l0bl8 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b8c609 l0bl8 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b8c610 l0bl8 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b8c611 l0bl8 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b8c612 l0bl8 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b8c613 l0bl8 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b8c614 l0bl8 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b8c615 l0bl8 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b8c616 l0bl8 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b8c617 l0bl8 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b8c618 l0bl8 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b8c619 l0bl8 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b8c620 l0bl8 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b8c621 l0bl8 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b8c622 l0bl8 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b8c623 l0bl8 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b8c624 l0bl8 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b8c625 l0bl8 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b8c626 l0bl8 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b8c627 l0bl8 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b8c628 l0bl8 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b8c629 l0bl8 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b8c630 l0bl8 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b8c631 l0bl8 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b8c632 l0bl8 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b8c633 l0bl8 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b8c634 l0bl8 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b8c635 l0bl8 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b8c636 l0bl8 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b8c637 l0bl8 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b8c638 l0bl8 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b8c639 l0bl8 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b8c640 l0bl8 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b8c641 l0bl8 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b8c642 l0bl8 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b8c643 l0bl8 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b8c644 l0bl8 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b8c645 l0bl8 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b8c646 l0bl8 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b8c647 l0bl8 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b8c648 l0bl8 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b8c649 l0bl8 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b8c650 l0bl8 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b8c651 l0bl8 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b8c652 l0bl8 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b8c653 l0bl8 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b8c654 l0bl8 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b8c655 l0bl8 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b8c656 l0bl8 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b8c657 l0bl8 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b8c658 l0bl8 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b8c659 l0bl8 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b8c660 l0bl8 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b8c661 l0bl8 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b8c662 l0bl8 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b8c663 l0bl8 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b8c664 l0bl8 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b8c665 l0bl8 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b8c666 l0bl8 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b8c667 l0bl8 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b8c668 l0bl8 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b8c669 l0bl8 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b8c670 l0bl8 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b8c671 l0bl8 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b8c672 l0bl8 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b8c673 l0bl8 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b8c674 l0bl8 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b8c675 l0bl8 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b8c676 l0bl8 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b8c677 l0bl8 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b8c678 l0bl8 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b8c679 l0bl8 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b8c680 l0bl8 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b8c681 l0bl8 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b8c682 l0bl8 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b8c683 l0bl8 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b8c684 l0bl8 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b8c685 l0bl8 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b8c686 l0bl8 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b8c687 l0bl8 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b8c688 l0bl8 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b8c689 l0bl8 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b8c690 l0bl8 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b8c691 l0bl8 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b8c692 l0bl8 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b8c693 l0bl8 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b8c694 l0bl8 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b8c695 l0bl8 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b8c696 l0bl8 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b8c697 l0bl8 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b8c698 l0bl8 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b8c699 l0bl8 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b8c700 l0bl8 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b8c701 l0bl8 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b8c702 l0bl8 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b8c703 l0bl8 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b8c704 l0bl8 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b8c705 l0bl8 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b8c706 l0bl8 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b8c707 l0bl8 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b8c708 l0bl8 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b8c709 l0bl8 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b8c710 l0bl8 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b8c711 l0bl8 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b8c712 l0bl8 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b8c713 l0bl8 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b8c714 l0bl8 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b8c715 l0bl8 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b8c716 l0bl8 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b8c717 l0bl8 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b8c718 l0bl8 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b8c719 l0bl8 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b8c720 l0bl8 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b8c721 l0bl8 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b8c722 l0bl8 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b8c723 l0bl8 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b8c724 l0bl8 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b8c725 l0bl8 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b8c726 l0bl8 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b8c727 l0bl8 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b8c728 l0bl8 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b8c729 l0bl8 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b8c730 l0bl8 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b8c731 l0bl8 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b8c732 l0bl8 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b8c733 l0bl8 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b8c734 l0bl8 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b8c735 l0bl8 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b8c736 l0bl8 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b8c737 l0bl8 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b8c738 l0bl8 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b8c739 l0bl8 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b8c740 l0bl8 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b8c741 l0bl8 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b8c742 l0bl8 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b8c743 l0bl8 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b8c744 l0bl8 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b8c745 l0bl8 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b8c746 l0bl8 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b8c747 l0bl8 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b8c748 l0bl8 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b8c749 l0bl8 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b8c750 l0bl8 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b8c751 l0bl8 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b8c752 l0bl8 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b8c753 l0bl8 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b8c754 l0bl8 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b8c755 l0bl8 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b8c756 l0bl8 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b8c757 l0bl8 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b8c758 l0bl8 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b8c759 l0bl8 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b8c760 l0bl8 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b8c761 l0bl8 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b8c762 l0bl8 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b8c763 l0bl8 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b8c764 l0bl8 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b8c765 l0bl8 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b8c766 l0bl8 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b8c767 l0bl8 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b8c768 l0bl8 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b8c769 l0bl8 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b8c770 l0bl8 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b8c771 l0bl8 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b8c772 l0bl8 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b8c773 l0bl8 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b8c774 l0bl8 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b8c775 l0bl8 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b8c776 l0bl8 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b8c777 l0bl8 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b8c778 l0bl8 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b8c779 l0bl8 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b8c780 l0bl8 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b8c781 l0bl8 vdd x781 x781b CELLD r1=10000e3 r0=900e3
xl0b8c782 l0bl8 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b8c783 l0bl8 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b9c0 l0bl9 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b9c1 l0bl9 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b9c2 l0bl9 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b9c3 l0bl9 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b9c4 l0bl9 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b9c5 l0bl9 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b9c6 l0bl9 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b9c7 l0bl9 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b9c8 l0bl9 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b9c9 l0bl9 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b9c10 l0bl9 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b9c11 l0bl9 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b9c12 l0bl9 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b9c13 l0bl9 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b9c14 l0bl9 vdd x14 x14b CELLD r1=10000e3 r0=900e3
xl0b9c15 l0bl9 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b9c16 l0bl9 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b9c17 l0bl9 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b9c18 l0bl9 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b9c19 l0bl9 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b9c20 l0bl9 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b9c21 l0bl9 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b9c22 l0bl9 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b9c23 l0bl9 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b9c24 l0bl9 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b9c25 l0bl9 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b9c26 l0bl9 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b9c27 l0bl9 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b9c28 l0bl9 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b9c29 l0bl9 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b9c30 l0bl9 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b9c31 l0bl9 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b9c32 l0bl9 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b9c33 l0bl9 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b9c34 l0bl9 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b9c35 l0bl9 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b9c36 l0bl9 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b9c37 l0bl9 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b9c38 l0bl9 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b9c39 l0bl9 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b9c40 l0bl9 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b9c41 l0bl9 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b9c42 l0bl9 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b9c43 l0bl9 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b9c44 l0bl9 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b9c45 l0bl9 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b9c46 l0bl9 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b9c47 l0bl9 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b9c48 l0bl9 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b9c49 l0bl9 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b9c50 l0bl9 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b9c51 l0bl9 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b9c52 l0bl9 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b9c53 l0bl9 vdd x53 x53b CELLD r1=900e3 r0=10000e3
xl0b9c54 l0bl9 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b9c55 l0bl9 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b9c56 l0bl9 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b9c57 l0bl9 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b9c58 l0bl9 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b9c59 l0bl9 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b9c60 l0bl9 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b9c61 l0bl9 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b9c62 l0bl9 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b9c63 l0bl9 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b9c64 l0bl9 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b9c65 l0bl9 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b9c66 l0bl9 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b9c67 l0bl9 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b9c68 l0bl9 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b9c69 l0bl9 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b9c70 l0bl9 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b9c71 l0bl9 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b9c72 l0bl9 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b9c73 l0bl9 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b9c74 l0bl9 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b9c75 l0bl9 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b9c76 l0bl9 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b9c77 l0bl9 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b9c78 l0bl9 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b9c79 l0bl9 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b9c80 l0bl9 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b9c81 l0bl9 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b9c82 l0bl9 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b9c83 l0bl9 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b9c84 l0bl9 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b9c85 l0bl9 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b9c86 l0bl9 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b9c87 l0bl9 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b9c88 l0bl9 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b9c89 l0bl9 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b9c90 l0bl9 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b9c91 l0bl9 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b9c92 l0bl9 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b9c93 l0bl9 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b9c94 l0bl9 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b9c95 l0bl9 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b9c96 l0bl9 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b9c97 l0bl9 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b9c98 l0bl9 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b9c99 l0bl9 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b9c100 l0bl9 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b9c101 l0bl9 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b9c102 l0bl9 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b9c103 l0bl9 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b9c104 l0bl9 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b9c105 l0bl9 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b9c106 l0bl9 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b9c107 l0bl9 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b9c108 l0bl9 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b9c109 l0bl9 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b9c110 l0bl9 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b9c111 l0bl9 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b9c112 l0bl9 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b9c113 l0bl9 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b9c114 l0bl9 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b9c115 l0bl9 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b9c116 l0bl9 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b9c117 l0bl9 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b9c118 l0bl9 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b9c119 l0bl9 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b9c120 l0bl9 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b9c121 l0bl9 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b9c122 l0bl9 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b9c123 l0bl9 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b9c124 l0bl9 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b9c125 l0bl9 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b9c126 l0bl9 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b9c127 l0bl9 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b9c128 l0bl9 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b9c129 l0bl9 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b9c130 l0bl9 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b9c131 l0bl9 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b9c132 l0bl9 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b9c133 l0bl9 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b9c134 l0bl9 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b9c135 l0bl9 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b9c136 l0bl9 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b9c137 l0bl9 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b9c138 l0bl9 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b9c139 l0bl9 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b9c140 l0bl9 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b9c141 l0bl9 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b9c142 l0bl9 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b9c143 l0bl9 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b9c144 l0bl9 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b9c145 l0bl9 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b9c146 l0bl9 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b9c147 l0bl9 vdd x147 x147b CELLD r1=900e3 r0=10000e3
xl0b9c148 l0bl9 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b9c149 l0bl9 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b9c150 l0bl9 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b9c151 l0bl9 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b9c152 l0bl9 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b9c153 l0bl9 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b9c154 l0bl9 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b9c155 l0bl9 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b9c156 l0bl9 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b9c157 l0bl9 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b9c158 l0bl9 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b9c159 l0bl9 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b9c160 l0bl9 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b9c161 l0bl9 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b9c162 l0bl9 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b9c163 l0bl9 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b9c164 l0bl9 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b9c165 l0bl9 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b9c166 l0bl9 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b9c167 l0bl9 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b9c168 l0bl9 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b9c169 l0bl9 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b9c170 l0bl9 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b9c171 l0bl9 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b9c172 l0bl9 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b9c173 l0bl9 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b9c174 l0bl9 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b9c175 l0bl9 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b9c176 l0bl9 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b9c177 l0bl9 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b9c178 l0bl9 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b9c179 l0bl9 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b9c180 l0bl9 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b9c181 l0bl9 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b9c182 l0bl9 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b9c183 l0bl9 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b9c184 l0bl9 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b9c185 l0bl9 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b9c186 l0bl9 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b9c187 l0bl9 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b9c188 l0bl9 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b9c189 l0bl9 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b9c190 l0bl9 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b9c191 l0bl9 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b9c192 l0bl9 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b9c193 l0bl9 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b9c194 l0bl9 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b9c195 l0bl9 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b9c196 l0bl9 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b9c197 l0bl9 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b9c198 l0bl9 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b9c199 l0bl9 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b9c200 l0bl9 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b9c201 l0bl9 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b9c202 l0bl9 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b9c203 l0bl9 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b9c204 l0bl9 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b9c205 l0bl9 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b9c206 l0bl9 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b9c207 l0bl9 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b9c208 l0bl9 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b9c209 l0bl9 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b9c210 l0bl9 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b9c211 l0bl9 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b9c212 l0bl9 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b9c213 l0bl9 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b9c214 l0bl9 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b9c215 l0bl9 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b9c216 l0bl9 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b9c217 l0bl9 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b9c218 l0bl9 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b9c219 l0bl9 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b9c220 l0bl9 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b9c221 l0bl9 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b9c222 l0bl9 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b9c223 l0bl9 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b9c224 l0bl9 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b9c225 l0bl9 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b9c226 l0bl9 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b9c227 l0bl9 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b9c228 l0bl9 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b9c229 l0bl9 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b9c230 l0bl9 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b9c231 l0bl9 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b9c232 l0bl9 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b9c233 l0bl9 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b9c234 l0bl9 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b9c235 l0bl9 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b9c236 l0bl9 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b9c237 l0bl9 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b9c238 l0bl9 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b9c239 l0bl9 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b9c240 l0bl9 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b9c241 l0bl9 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b9c242 l0bl9 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b9c243 l0bl9 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b9c244 l0bl9 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b9c245 l0bl9 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b9c246 l0bl9 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b9c247 l0bl9 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b9c248 l0bl9 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b9c249 l0bl9 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b9c250 l0bl9 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b9c251 l0bl9 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b9c252 l0bl9 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b9c253 l0bl9 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b9c254 l0bl9 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b9c255 l0bl9 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b9c256 l0bl9 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b9c257 l0bl9 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b9c258 l0bl9 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b9c259 l0bl9 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b9c260 l0bl9 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b9c261 l0bl9 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b9c262 l0bl9 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b9c263 l0bl9 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b9c264 l0bl9 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b9c265 l0bl9 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b9c266 l0bl9 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b9c267 l0bl9 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b9c268 l0bl9 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b9c269 l0bl9 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b9c270 l0bl9 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b9c271 l0bl9 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b9c272 l0bl9 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b9c273 l0bl9 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b9c274 l0bl9 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b9c275 l0bl9 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b9c276 l0bl9 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b9c277 l0bl9 vdd x277 x277b CELLD r1=900e3 r0=10000e3
xl0b9c278 l0bl9 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b9c279 l0bl9 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b9c280 l0bl9 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b9c281 l0bl9 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b9c282 l0bl9 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b9c283 l0bl9 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b9c284 l0bl9 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b9c285 l0bl9 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b9c286 l0bl9 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b9c287 l0bl9 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b9c288 l0bl9 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b9c289 l0bl9 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b9c290 l0bl9 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b9c291 l0bl9 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b9c292 l0bl9 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b9c293 l0bl9 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b9c294 l0bl9 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b9c295 l0bl9 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b9c296 l0bl9 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b9c297 l0bl9 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b9c298 l0bl9 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b9c299 l0bl9 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b9c300 l0bl9 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b9c301 l0bl9 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b9c302 l0bl9 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b9c303 l0bl9 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b9c304 l0bl9 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b9c305 l0bl9 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b9c306 l0bl9 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b9c307 l0bl9 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b9c308 l0bl9 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b9c309 l0bl9 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b9c310 l0bl9 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b9c311 l0bl9 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b9c312 l0bl9 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b9c313 l0bl9 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b9c314 l0bl9 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b9c315 l0bl9 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b9c316 l0bl9 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b9c317 l0bl9 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b9c318 l0bl9 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b9c319 l0bl9 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b9c320 l0bl9 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b9c321 l0bl9 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b9c322 l0bl9 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b9c323 l0bl9 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b9c324 l0bl9 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b9c325 l0bl9 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b9c326 l0bl9 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b9c327 l0bl9 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b9c328 l0bl9 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b9c329 l0bl9 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b9c330 l0bl9 vdd x330 x330b CELLD r1=900e3 r0=10000e3
xl0b9c331 l0bl9 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b9c332 l0bl9 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b9c333 l0bl9 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b9c334 l0bl9 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b9c335 l0bl9 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b9c336 l0bl9 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b9c337 l0bl9 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b9c338 l0bl9 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b9c339 l0bl9 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b9c340 l0bl9 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b9c341 l0bl9 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b9c342 l0bl9 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b9c343 l0bl9 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b9c344 l0bl9 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b9c345 l0bl9 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b9c346 l0bl9 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b9c347 l0bl9 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b9c348 l0bl9 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b9c349 l0bl9 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b9c350 l0bl9 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b9c351 l0bl9 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b9c352 l0bl9 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b9c353 l0bl9 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b9c354 l0bl9 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b9c355 l0bl9 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b9c356 l0bl9 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b9c357 l0bl9 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b9c358 l0bl9 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b9c359 l0bl9 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b9c360 l0bl9 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b9c361 l0bl9 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b9c362 l0bl9 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b9c363 l0bl9 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b9c364 l0bl9 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b9c365 l0bl9 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b9c366 l0bl9 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b9c367 l0bl9 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b9c368 l0bl9 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b9c369 l0bl9 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b9c370 l0bl9 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b9c371 l0bl9 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b9c372 l0bl9 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b9c373 l0bl9 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b9c374 l0bl9 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b9c375 l0bl9 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b9c376 l0bl9 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b9c377 l0bl9 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b9c378 l0bl9 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b9c379 l0bl9 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b9c380 l0bl9 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b9c381 l0bl9 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b9c382 l0bl9 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b9c383 l0bl9 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b9c384 l0bl9 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b9c385 l0bl9 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b9c386 l0bl9 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b9c387 l0bl9 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b9c388 l0bl9 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b9c389 l0bl9 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b9c390 l0bl9 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b9c391 l0bl9 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b9c392 l0bl9 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b9c393 l0bl9 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b9c394 l0bl9 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b9c395 l0bl9 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b9c396 l0bl9 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b9c397 l0bl9 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b9c398 l0bl9 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b9c399 l0bl9 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b9c400 l0bl9 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b9c401 l0bl9 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b9c402 l0bl9 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b9c403 l0bl9 vdd x403 x403b CELLD r1=10000e3 r0=900e3
xl0b9c404 l0bl9 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b9c405 l0bl9 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b9c406 l0bl9 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b9c407 l0bl9 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b9c408 l0bl9 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b9c409 l0bl9 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b9c410 l0bl9 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b9c411 l0bl9 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b9c412 l0bl9 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b9c413 l0bl9 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b9c414 l0bl9 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b9c415 l0bl9 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b9c416 l0bl9 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b9c417 l0bl9 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b9c418 l0bl9 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b9c419 l0bl9 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b9c420 l0bl9 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b9c421 l0bl9 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b9c422 l0bl9 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b9c423 l0bl9 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b9c424 l0bl9 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b9c425 l0bl9 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b9c426 l0bl9 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b9c427 l0bl9 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b9c428 l0bl9 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b9c429 l0bl9 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b9c430 l0bl9 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b9c431 l0bl9 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b9c432 l0bl9 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b9c433 l0bl9 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b9c434 l0bl9 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b9c435 l0bl9 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b9c436 l0bl9 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b9c437 l0bl9 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b9c438 l0bl9 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b9c439 l0bl9 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b9c440 l0bl9 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b9c441 l0bl9 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b9c442 l0bl9 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b9c443 l0bl9 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b9c444 l0bl9 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b9c445 l0bl9 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b9c446 l0bl9 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b9c447 l0bl9 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b9c448 l0bl9 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b9c449 l0bl9 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b9c450 l0bl9 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b9c451 l0bl9 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b9c452 l0bl9 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b9c453 l0bl9 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b9c454 l0bl9 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b9c455 l0bl9 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b9c456 l0bl9 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b9c457 l0bl9 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b9c458 l0bl9 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b9c459 l0bl9 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b9c460 l0bl9 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b9c461 l0bl9 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b9c462 l0bl9 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b9c463 l0bl9 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b9c464 l0bl9 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b9c465 l0bl9 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b9c466 l0bl9 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b9c467 l0bl9 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b9c468 l0bl9 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b9c469 l0bl9 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b9c470 l0bl9 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b9c471 l0bl9 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b9c472 l0bl9 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b9c473 l0bl9 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b9c474 l0bl9 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b9c475 l0bl9 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b9c476 l0bl9 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b9c477 l0bl9 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b9c478 l0bl9 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b9c479 l0bl9 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b9c480 l0bl9 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b9c481 l0bl9 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b9c482 l0bl9 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b9c483 l0bl9 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b9c484 l0bl9 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b9c485 l0bl9 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b9c486 l0bl9 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b9c487 l0bl9 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b9c488 l0bl9 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b9c489 l0bl9 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b9c490 l0bl9 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b9c491 l0bl9 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b9c492 l0bl9 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b9c493 l0bl9 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b9c494 l0bl9 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b9c495 l0bl9 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b9c496 l0bl9 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b9c497 l0bl9 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b9c498 l0bl9 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b9c499 l0bl9 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b9c500 l0bl9 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b9c501 l0bl9 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b9c502 l0bl9 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b9c503 l0bl9 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b9c504 l0bl9 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b9c505 l0bl9 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b9c506 l0bl9 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b9c507 l0bl9 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b9c508 l0bl9 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b9c509 l0bl9 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b9c510 l0bl9 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b9c511 l0bl9 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b9c512 l0bl9 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b9c513 l0bl9 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b9c514 l0bl9 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b9c515 l0bl9 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b9c516 l0bl9 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b9c517 l0bl9 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b9c518 l0bl9 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b9c519 l0bl9 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b9c520 l0bl9 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b9c521 l0bl9 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b9c522 l0bl9 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b9c523 l0bl9 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b9c524 l0bl9 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b9c525 l0bl9 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b9c526 l0bl9 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b9c527 l0bl9 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b9c528 l0bl9 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b9c529 l0bl9 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b9c530 l0bl9 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b9c531 l0bl9 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b9c532 l0bl9 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b9c533 l0bl9 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b9c534 l0bl9 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b9c535 l0bl9 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b9c536 l0bl9 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b9c537 l0bl9 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b9c538 l0bl9 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b9c539 l0bl9 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b9c540 l0bl9 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b9c541 l0bl9 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b9c542 l0bl9 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b9c543 l0bl9 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b9c544 l0bl9 vdd x544 x544b CELLD r1=10000e3 r0=900e3
xl0b9c545 l0bl9 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b9c546 l0bl9 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b9c547 l0bl9 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b9c548 l0bl9 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b9c549 l0bl9 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b9c550 l0bl9 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b9c551 l0bl9 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b9c552 l0bl9 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b9c553 l0bl9 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b9c554 l0bl9 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b9c555 l0bl9 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b9c556 l0bl9 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b9c557 l0bl9 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b9c558 l0bl9 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b9c559 l0bl9 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b9c560 l0bl9 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b9c561 l0bl9 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b9c562 l0bl9 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b9c563 l0bl9 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b9c564 l0bl9 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b9c565 l0bl9 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b9c566 l0bl9 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b9c567 l0bl9 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b9c568 l0bl9 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b9c569 l0bl9 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b9c570 l0bl9 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b9c571 l0bl9 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b9c572 l0bl9 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b9c573 l0bl9 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b9c574 l0bl9 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b9c575 l0bl9 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b9c576 l0bl9 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b9c577 l0bl9 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b9c578 l0bl9 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b9c579 l0bl9 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b9c580 l0bl9 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b9c581 l0bl9 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b9c582 l0bl9 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b9c583 l0bl9 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b9c584 l0bl9 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b9c585 l0bl9 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b9c586 l0bl9 vdd x586 x586b CELLD r1=10000e3 r0=900e3
xl0b9c587 l0bl9 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b9c588 l0bl9 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b9c589 l0bl9 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b9c590 l0bl9 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b9c591 l0bl9 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b9c592 l0bl9 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b9c593 l0bl9 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b9c594 l0bl9 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b9c595 l0bl9 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b9c596 l0bl9 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b9c597 l0bl9 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b9c598 l0bl9 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b9c599 l0bl9 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b9c600 l0bl9 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b9c601 l0bl9 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b9c602 l0bl9 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b9c603 l0bl9 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b9c604 l0bl9 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b9c605 l0bl9 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b9c606 l0bl9 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b9c607 l0bl9 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b9c608 l0bl9 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b9c609 l0bl9 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b9c610 l0bl9 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b9c611 l0bl9 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b9c612 l0bl9 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b9c613 l0bl9 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b9c614 l0bl9 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b9c615 l0bl9 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b9c616 l0bl9 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b9c617 l0bl9 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b9c618 l0bl9 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b9c619 l0bl9 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b9c620 l0bl9 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b9c621 l0bl9 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b9c622 l0bl9 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b9c623 l0bl9 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b9c624 l0bl9 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b9c625 l0bl9 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b9c626 l0bl9 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b9c627 l0bl9 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b9c628 l0bl9 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b9c629 l0bl9 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b9c630 l0bl9 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b9c631 l0bl9 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b9c632 l0bl9 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b9c633 l0bl9 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b9c634 l0bl9 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b9c635 l0bl9 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b9c636 l0bl9 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b9c637 l0bl9 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b9c638 l0bl9 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b9c639 l0bl9 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b9c640 l0bl9 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b9c641 l0bl9 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b9c642 l0bl9 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b9c643 l0bl9 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b9c644 l0bl9 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b9c645 l0bl9 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b9c646 l0bl9 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b9c647 l0bl9 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b9c648 l0bl9 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b9c649 l0bl9 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b9c650 l0bl9 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b9c651 l0bl9 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b9c652 l0bl9 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b9c653 l0bl9 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b9c654 l0bl9 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b9c655 l0bl9 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b9c656 l0bl9 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b9c657 l0bl9 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b9c658 l0bl9 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b9c659 l0bl9 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b9c660 l0bl9 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b9c661 l0bl9 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b9c662 l0bl9 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b9c663 l0bl9 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b9c664 l0bl9 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b9c665 l0bl9 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b9c666 l0bl9 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b9c667 l0bl9 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b9c668 l0bl9 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b9c669 l0bl9 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b9c670 l0bl9 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b9c671 l0bl9 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b9c672 l0bl9 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b9c673 l0bl9 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b9c674 l0bl9 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b9c675 l0bl9 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b9c676 l0bl9 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b9c677 l0bl9 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b9c678 l0bl9 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b9c679 l0bl9 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b9c680 l0bl9 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b9c681 l0bl9 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b9c682 l0bl9 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b9c683 l0bl9 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b9c684 l0bl9 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b9c685 l0bl9 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b9c686 l0bl9 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b9c687 l0bl9 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b9c688 l0bl9 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b9c689 l0bl9 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b9c690 l0bl9 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b9c691 l0bl9 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b9c692 l0bl9 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b9c693 l0bl9 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b9c694 l0bl9 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b9c695 l0bl9 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b9c696 l0bl9 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b9c697 l0bl9 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b9c698 l0bl9 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b9c699 l0bl9 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b9c700 l0bl9 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b9c701 l0bl9 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b9c702 l0bl9 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b9c703 l0bl9 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b9c704 l0bl9 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b9c705 l0bl9 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b9c706 l0bl9 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b9c707 l0bl9 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b9c708 l0bl9 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b9c709 l0bl9 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b9c710 l0bl9 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b9c711 l0bl9 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b9c712 l0bl9 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b9c713 l0bl9 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b9c714 l0bl9 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b9c715 l0bl9 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b9c716 l0bl9 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b9c717 l0bl9 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b9c718 l0bl9 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b9c719 l0bl9 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b9c720 l0bl9 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b9c721 l0bl9 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b9c722 l0bl9 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b9c723 l0bl9 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b9c724 l0bl9 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b9c725 l0bl9 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b9c726 l0bl9 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b9c727 l0bl9 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b9c728 l0bl9 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b9c729 l0bl9 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b9c730 l0bl9 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b9c731 l0bl9 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b9c732 l0bl9 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b9c733 l0bl9 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b9c734 l0bl9 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b9c735 l0bl9 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b9c736 l0bl9 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b9c737 l0bl9 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b9c738 l0bl9 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b9c739 l0bl9 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b9c740 l0bl9 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b9c741 l0bl9 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b9c742 l0bl9 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b9c743 l0bl9 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b9c744 l0bl9 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b9c745 l0bl9 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b9c746 l0bl9 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b9c747 l0bl9 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b9c748 l0bl9 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b9c749 l0bl9 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b9c750 l0bl9 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b9c751 l0bl9 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b9c752 l0bl9 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b9c753 l0bl9 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b9c754 l0bl9 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b9c755 l0bl9 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b9c756 l0bl9 vdd x756 x756b CELLD r1=900e3 r0=10000e3
xl0b9c757 l0bl9 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b9c758 l0bl9 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b9c759 l0bl9 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b9c760 l0bl9 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b9c761 l0bl9 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b9c762 l0bl9 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b9c763 l0bl9 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b9c764 l0bl9 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b9c765 l0bl9 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b9c766 l0bl9 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b9c767 l0bl9 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b9c768 l0bl9 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b9c769 l0bl9 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b9c770 l0bl9 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b9c771 l0bl9 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b9c772 l0bl9 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b9c773 l0bl9 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b9c774 l0bl9 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b9c775 l0bl9 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b9c776 l0bl9 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b9c777 l0bl9 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b9c778 l0bl9 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b9c779 l0bl9 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b9c780 l0bl9 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b9c781 l0bl9 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b9c782 l0bl9 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b9c783 l0bl9 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b10c0 l0bl10 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b10c1 l0bl10 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b10c2 l0bl10 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b10c3 l0bl10 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b10c4 l0bl10 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b10c5 l0bl10 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b10c6 l0bl10 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b10c7 l0bl10 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b10c8 l0bl10 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b10c9 l0bl10 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b10c10 l0bl10 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b10c11 l0bl10 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b10c12 l0bl10 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b10c13 l0bl10 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b10c14 l0bl10 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b10c15 l0bl10 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b10c16 l0bl10 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b10c17 l0bl10 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b10c18 l0bl10 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b10c19 l0bl10 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b10c20 l0bl10 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b10c21 l0bl10 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b10c22 l0bl10 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b10c23 l0bl10 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b10c24 l0bl10 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b10c25 l0bl10 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b10c26 l0bl10 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b10c27 l0bl10 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b10c28 l0bl10 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b10c29 l0bl10 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b10c30 l0bl10 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b10c31 l0bl10 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b10c32 l0bl10 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b10c33 l0bl10 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b10c34 l0bl10 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b10c35 l0bl10 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b10c36 l0bl10 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b10c37 l0bl10 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b10c38 l0bl10 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b10c39 l0bl10 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b10c40 l0bl10 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b10c41 l0bl10 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b10c42 l0bl10 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b10c43 l0bl10 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b10c44 l0bl10 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b10c45 l0bl10 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b10c46 l0bl10 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b10c47 l0bl10 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b10c48 l0bl10 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b10c49 l0bl10 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b10c50 l0bl10 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b10c51 l0bl10 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b10c52 l0bl10 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b10c53 l0bl10 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b10c54 l0bl10 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b10c55 l0bl10 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b10c56 l0bl10 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b10c57 l0bl10 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b10c58 l0bl10 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b10c59 l0bl10 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b10c60 l0bl10 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b10c61 l0bl10 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b10c62 l0bl10 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b10c63 l0bl10 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b10c64 l0bl10 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b10c65 l0bl10 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b10c66 l0bl10 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b10c67 l0bl10 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b10c68 l0bl10 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b10c69 l0bl10 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b10c70 l0bl10 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b10c71 l0bl10 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b10c72 l0bl10 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b10c73 l0bl10 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b10c74 l0bl10 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b10c75 l0bl10 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b10c76 l0bl10 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b10c77 l0bl10 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b10c78 l0bl10 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b10c79 l0bl10 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b10c80 l0bl10 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b10c81 l0bl10 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b10c82 l0bl10 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b10c83 l0bl10 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b10c84 l0bl10 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b10c85 l0bl10 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b10c86 l0bl10 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b10c87 l0bl10 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b10c88 l0bl10 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b10c89 l0bl10 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b10c90 l0bl10 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b10c91 l0bl10 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b10c92 l0bl10 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b10c93 l0bl10 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b10c94 l0bl10 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b10c95 l0bl10 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b10c96 l0bl10 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b10c97 l0bl10 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b10c98 l0bl10 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b10c99 l0bl10 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b10c100 l0bl10 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b10c101 l0bl10 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b10c102 l0bl10 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b10c103 l0bl10 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b10c104 l0bl10 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b10c105 l0bl10 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b10c106 l0bl10 vdd x106 x106b CELLD r1=10000e3 r0=900e3
xl0b10c107 l0bl10 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b10c108 l0bl10 vdd x108 x108b CELLD r1=10000e3 r0=900e3
xl0b10c109 l0bl10 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b10c110 l0bl10 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b10c111 l0bl10 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b10c112 l0bl10 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b10c113 l0bl10 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b10c114 l0bl10 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b10c115 l0bl10 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b10c116 l0bl10 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b10c117 l0bl10 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b10c118 l0bl10 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b10c119 l0bl10 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b10c120 l0bl10 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b10c121 l0bl10 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b10c122 l0bl10 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b10c123 l0bl10 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b10c124 l0bl10 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b10c125 l0bl10 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b10c126 l0bl10 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b10c127 l0bl10 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b10c128 l0bl10 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b10c129 l0bl10 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b10c130 l0bl10 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b10c131 l0bl10 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b10c132 l0bl10 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b10c133 l0bl10 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b10c134 l0bl10 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b10c135 l0bl10 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b10c136 l0bl10 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b10c137 l0bl10 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b10c138 l0bl10 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b10c139 l0bl10 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b10c140 l0bl10 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b10c141 l0bl10 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b10c142 l0bl10 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b10c143 l0bl10 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b10c144 l0bl10 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b10c145 l0bl10 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b10c146 l0bl10 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b10c147 l0bl10 vdd x147 x147b CELLD r1=900e3 r0=10000e3
xl0b10c148 l0bl10 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b10c149 l0bl10 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b10c150 l0bl10 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b10c151 l0bl10 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b10c152 l0bl10 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b10c153 l0bl10 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b10c154 l0bl10 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b10c155 l0bl10 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b10c156 l0bl10 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b10c157 l0bl10 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b10c158 l0bl10 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b10c159 l0bl10 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b10c160 l0bl10 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b10c161 l0bl10 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b10c162 l0bl10 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b10c163 l0bl10 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b10c164 l0bl10 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b10c165 l0bl10 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b10c166 l0bl10 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b10c167 l0bl10 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b10c168 l0bl10 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b10c169 l0bl10 vdd x169 x169b CELLD r1=10000e3 r0=900e3
xl0b10c170 l0bl10 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b10c171 l0bl10 vdd x171 x171b CELLD r1=10000e3 r0=900e3
xl0b10c172 l0bl10 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b10c173 l0bl10 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b10c174 l0bl10 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b10c175 l0bl10 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b10c176 l0bl10 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b10c177 l0bl10 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b10c178 l0bl10 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b10c179 l0bl10 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b10c180 l0bl10 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b10c181 l0bl10 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b10c182 l0bl10 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b10c183 l0bl10 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b10c184 l0bl10 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b10c185 l0bl10 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b10c186 l0bl10 vdd x186 x186b CELLD r1=10000e3 r0=900e3
xl0b10c187 l0bl10 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b10c188 l0bl10 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b10c189 l0bl10 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b10c190 l0bl10 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b10c191 l0bl10 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b10c192 l0bl10 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b10c193 l0bl10 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b10c194 l0bl10 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b10c195 l0bl10 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b10c196 l0bl10 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b10c197 l0bl10 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b10c198 l0bl10 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b10c199 l0bl10 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b10c200 l0bl10 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b10c201 l0bl10 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b10c202 l0bl10 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b10c203 l0bl10 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b10c204 l0bl10 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b10c205 l0bl10 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b10c206 l0bl10 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b10c207 l0bl10 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b10c208 l0bl10 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b10c209 l0bl10 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b10c210 l0bl10 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b10c211 l0bl10 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b10c212 l0bl10 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b10c213 l0bl10 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b10c214 l0bl10 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b10c215 l0bl10 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b10c216 l0bl10 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b10c217 l0bl10 vdd x217 x217b CELLD r1=900e3 r0=10000e3
xl0b10c218 l0bl10 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b10c219 l0bl10 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b10c220 l0bl10 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b10c221 l0bl10 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b10c222 l0bl10 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b10c223 l0bl10 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b10c224 l0bl10 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b10c225 l0bl10 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b10c226 l0bl10 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b10c227 l0bl10 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b10c228 l0bl10 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b10c229 l0bl10 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b10c230 l0bl10 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b10c231 l0bl10 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b10c232 l0bl10 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b10c233 l0bl10 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b10c234 l0bl10 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b10c235 l0bl10 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b10c236 l0bl10 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b10c237 l0bl10 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b10c238 l0bl10 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b10c239 l0bl10 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b10c240 l0bl10 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b10c241 l0bl10 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b10c242 l0bl10 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b10c243 l0bl10 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b10c244 l0bl10 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b10c245 l0bl10 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b10c246 l0bl10 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b10c247 l0bl10 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b10c248 l0bl10 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b10c249 l0bl10 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b10c250 l0bl10 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b10c251 l0bl10 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b10c252 l0bl10 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b10c253 l0bl10 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b10c254 l0bl10 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b10c255 l0bl10 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b10c256 l0bl10 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b10c257 l0bl10 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b10c258 l0bl10 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b10c259 l0bl10 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b10c260 l0bl10 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b10c261 l0bl10 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b10c262 l0bl10 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b10c263 l0bl10 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b10c264 l0bl10 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b10c265 l0bl10 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b10c266 l0bl10 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b10c267 l0bl10 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b10c268 l0bl10 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b10c269 l0bl10 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b10c270 l0bl10 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b10c271 l0bl10 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b10c272 l0bl10 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b10c273 l0bl10 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b10c274 l0bl10 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b10c275 l0bl10 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b10c276 l0bl10 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b10c277 l0bl10 vdd x277 x277b CELLD r1=900e3 r0=10000e3
xl0b10c278 l0bl10 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b10c279 l0bl10 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b10c280 l0bl10 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b10c281 l0bl10 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b10c282 l0bl10 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b10c283 l0bl10 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b10c284 l0bl10 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b10c285 l0bl10 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b10c286 l0bl10 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b10c287 l0bl10 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b10c288 l0bl10 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b10c289 l0bl10 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b10c290 l0bl10 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b10c291 l0bl10 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b10c292 l0bl10 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b10c293 l0bl10 vdd x293 x293b CELLD r1=900e3 r0=10000e3
xl0b10c294 l0bl10 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b10c295 l0bl10 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b10c296 l0bl10 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b10c297 l0bl10 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b10c298 l0bl10 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b10c299 l0bl10 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b10c300 l0bl10 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b10c301 l0bl10 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b10c302 l0bl10 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b10c303 l0bl10 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b10c304 l0bl10 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b10c305 l0bl10 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b10c306 l0bl10 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b10c307 l0bl10 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b10c308 l0bl10 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b10c309 l0bl10 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b10c310 l0bl10 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b10c311 l0bl10 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b10c312 l0bl10 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b10c313 l0bl10 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b10c314 l0bl10 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b10c315 l0bl10 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b10c316 l0bl10 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b10c317 l0bl10 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b10c318 l0bl10 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b10c319 l0bl10 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b10c320 l0bl10 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b10c321 l0bl10 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b10c322 l0bl10 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b10c323 l0bl10 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b10c324 l0bl10 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b10c325 l0bl10 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b10c326 l0bl10 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b10c327 l0bl10 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b10c328 l0bl10 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b10c329 l0bl10 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b10c330 l0bl10 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b10c331 l0bl10 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b10c332 l0bl10 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b10c333 l0bl10 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b10c334 l0bl10 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b10c335 l0bl10 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b10c336 l0bl10 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b10c337 l0bl10 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b10c338 l0bl10 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b10c339 l0bl10 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b10c340 l0bl10 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b10c341 l0bl10 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b10c342 l0bl10 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b10c343 l0bl10 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b10c344 l0bl10 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b10c345 l0bl10 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b10c346 l0bl10 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b10c347 l0bl10 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b10c348 l0bl10 vdd x348 x348b CELLD r1=10000e3 r0=900e3
xl0b10c349 l0bl10 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b10c350 l0bl10 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b10c351 l0bl10 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b10c352 l0bl10 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b10c353 l0bl10 vdd x353 x353b CELLD r1=10000e3 r0=900e3
xl0b10c354 l0bl10 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b10c355 l0bl10 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b10c356 l0bl10 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b10c357 l0bl10 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b10c358 l0bl10 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b10c359 l0bl10 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b10c360 l0bl10 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b10c361 l0bl10 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b10c362 l0bl10 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b10c363 l0bl10 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b10c364 l0bl10 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b10c365 l0bl10 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b10c366 l0bl10 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b10c367 l0bl10 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b10c368 l0bl10 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b10c369 l0bl10 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b10c370 l0bl10 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b10c371 l0bl10 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b10c372 l0bl10 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b10c373 l0bl10 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b10c374 l0bl10 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b10c375 l0bl10 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b10c376 l0bl10 vdd x376 x376b CELLD r1=10000e3 r0=900e3
xl0b10c377 l0bl10 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b10c378 l0bl10 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b10c379 l0bl10 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b10c380 l0bl10 vdd x380 x380b CELLD r1=10000e3 r0=900e3
xl0b10c381 l0bl10 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b10c382 l0bl10 vdd x382 x382b CELLD r1=10000e3 r0=900e3
xl0b10c383 l0bl10 vdd x383 x383b CELLD r1=10000e3 r0=900e3
xl0b10c384 l0bl10 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b10c385 l0bl10 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b10c386 l0bl10 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b10c387 l0bl10 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b10c388 l0bl10 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b10c389 l0bl10 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b10c390 l0bl10 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b10c391 l0bl10 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b10c392 l0bl10 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b10c393 l0bl10 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b10c394 l0bl10 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b10c395 l0bl10 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b10c396 l0bl10 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b10c397 l0bl10 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b10c398 l0bl10 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b10c399 l0bl10 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b10c400 l0bl10 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b10c401 l0bl10 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b10c402 l0bl10 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b10c403 l0bl10 vdd x403 x403b CELLD r1=10000e3 r0=900e3
xl0b10c404 l0bl10 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b10c405 l0bl10 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b10c406 l0bl10 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b10c407 l0bl10 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b10c408 l0bl10 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b10c409 l0bl10 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b10c410 l0bl10 vdd x410 x410b CELLD r1=10000e3 r0=900e3
xl0b10c411 l0bl10 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b10c412 l0bl10 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b10c413 l0bl10 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b10c414 l0bl10 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b10c415 l0bl10 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b10c416 l0bl10 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b10c417 l0bl10 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b10c418 l0bl10 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b10c419 l0bl10 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b10c420 l0bl10 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b10c421 l0bl10 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b10c422 l0bl10 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b10c423 l0bl10 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b10c424 l0bl10 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b10c425 l0bl10 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b10c426 l0bl10 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b10c427 l0bl10 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b10c428 l0bl10 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b10c429 l0bl10 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b10c430 l0bl10 vdd x430 x430b CELLD r1=10000e3 r0=900e3
xl0b10c431 l0bl10 vdd x431 x431b CELLD r1=10000e3 r0=900e3
xl0b10c432 l0bl10 vdd x432 x432b CELLD r1=10000e3 r0=900e3
xl0b10c433 l0bl10 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b10c434 l0bl10 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b10c435 l0bl10 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b10c436 l0bl10 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b10c437 l0bl10 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b10c438 l0bl10 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b10c439 l0bl10 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b10c440 l0bl10 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b10c441 l0bl10 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b10c442 l0bl10 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b10c443 l0bl10 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b10c444 l0bl10 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b10c445 l0bl10 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b10c446 l0bl10 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b10c447 l0bl10 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b10c448 l0bl10 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b10c449 l0bl10 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b10c450 l0bl10 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b10c451 l0bl10 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b10c452 l0bl10 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b10c453 l0bl10 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b10c454 l0bl10 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b10c455 l0bl10 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b10c456 l0bl10 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b10c457 l0bl10 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b10c458 l0bl10 vdd x458 x458b CELLD r1=10000e3 r0=900e3
xl0b10c459 l0bl10 vdd x459 x459b CELLD r1=10000e3 r0=900e3
xl0b10c460 l0bl10 vdd x460 x460b CELLD r1=10000e3 r0=900e3
xl0b10c461 l0bl10 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b10c462 l0bl10 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b10c463 l0bl10 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b10c464 l0bl10 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b10c465 l0bl10 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b10c466 l0bl10 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b10c467 l0bl10 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b10c468 l0bl10 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b10c469 l0bl10 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b10c470 l0bl10 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b10c471 l0bl10 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b10c472 l0bl10 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b10c473 l0bl10 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b10c474 l0bl10 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b10c475 l0bl10 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b10c476 l0bl10 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b10c477 l0bl10 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b10c478 l0bl10 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b10c479 l0bl10 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b10c480 l0bl10 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b10c481 l0bl10 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b10c482 l0bl10 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b10c483 l0bl10 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b10c484 l0bl10 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b10c485 l0bl10 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b10c486 l0bl10 vdd x486 x486b CELLD r1=10000e3 r0=900e3
xl0b10c487 l0bl10 vdd x487 x487b CELLD r1=10000e3 r0=900e3
xl0b10c488 l0bl10 vdd x488 x488b CELLD r1=10000e3 r0=900e3
xl0b10c489 l0bl10 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b10c490 l0bl10 vdd x490 x490b CELLD r1=10000e3 r0=900e3
xl0b10c491 l0bl10 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b10c492 l0bl10 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b10c493 l0bl10 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b10c494 l0bl10 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b10c495 l0bl10 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b10c496 l0bl10 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b10c497 l0bl10 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b10c498 l0bl10 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b10c499 l0bl10 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b10c500 l0bl10 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b10c501 l0bl10 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b10c502 l0bl10 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b10c503 l0bl10 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b10c504 l0bl10 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b10c505 l0bl10 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b10c506 l0bl10 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b10c507 l0bl10 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b10c508 l0bl10 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b10c509 l0bl10 vdd x509 x509b CELLD r1=900e3 r0=10000e3
xl0b10c510 l0bl10 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b10c511 l0bl10 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b10c512 l0bl10 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b10c513 l0bl10 vdd x513 x513b CELLD r1=10000e3 r0=900e3
xl0b10c514 l0bl10 vdd x514 x514b CELLD r1=10000e3 r0=900e3
xl0b10c515 l0bl10 vdd x515 x515b CELLD r1=10000e3 r0=900e3
xl0b10c516 l0bl10 vdd x516 x516b CELLD r1=10000e3 r0=900e3
xl0b10c517 l0bl10 vdd x517 x517b CELLD r1=10000e3 r0=900e3
xl0b10c518 l0bl10 vdd x518 x518b CELLD r1=10000e3 r0=900e3
xl0b10c519 l0bl10 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b10c520 l0bl10 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b10c521 l0bl10 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b10c522 l0bl10 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b10c523 l0bl10 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b10c524 l0bl10 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b10c525 l0bl10 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b10c526 l0bl10 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b10c527 l0bl10 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b10c528 l0bl10 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b10c529 l0bl10 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b10c530 l0bl10 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b10c531 l0bl10 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b10c532 l0bl10 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b10c533 l0bl10 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b10c534 l0bl10 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b10c535 l0bl10 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b10c536 l0bl10 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b10c537 l0bl10 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b10c538 l0bl10 vdd x538 x538b CELLD r1=900e3 r0=10000e3
xl0b10c539 l0bl10 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b10c540 l0bl10 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b10c541 l0bl10 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b10c542 l0bl10 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b10c543 l0bl10 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b10c544 l0bl10 vdd x544 x544b CELLD r1=10000e3 r0=900e3
xl0b10c545 l0bl10 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b10c546 l0bl10 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b10c547 l0bl10 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b10c548 l0bl10 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b10c549 l0bl10 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b10c550 l0bl10 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b10c551 l0bl10 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b10c552 l0bl10 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b10c553 l0bl10 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b10c554 l0bl10 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b10c555 l0bl10 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b10c556 l0bl10 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b10c557 l0bl10 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b10c558 l0bl10 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b10c559 l0bl10 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b10c560 l0bl10 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b10c561 l0bl10 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b10c562 l0bl10 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b10c563 l0bl10 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b10c564 l0bl10 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b10c565 l0bl10 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b10c566 l0bl10 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b10c567 l0bl10 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b10c568 l0bl10 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b10c569 l0bl10 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b10c570 l0bl10 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b10c571 l0bl10 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b10c572 l0bl10 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b10c573 l0bl10 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b10c574 l0bl10 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b10c575 l0bl10 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b10c576 l0bl10 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b10c577 l0bl10 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b10c578 l0bl10 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b10c579 l0bl10 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b10c580 l0bl10 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b10c581 l0bl10 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b10c582 l0bl10 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b10c583 l0bl10 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b10c584 l0bl10 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b10c585 l0bl10 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b10c586 l0bl10 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b10c587 l0bl10 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b10c588 l0bl10 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b10c589 l0bl10 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b10c590 l0bl10 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b10c591 l0bl10 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b10c592 l0bl10 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b10c593 l0bl10 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b10c594 l0bl10 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b10c595 l0bl10 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b10c596 l0bl10 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b10c597 l0bl10 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b10c598 l0bl10 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b10c599 l0bl10 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b10c600 l0bl10 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b10c601 l0bl10 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b10c602 l0bl10 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b10c603 l0bl10 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b10c604 l0bl10 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b10c605 l0bl10 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b10c606 l0bl10 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b10c607 l0bl10 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b10c608 l0bl10 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b10c609 l0bl10 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b10c610 l0bl10 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b10c611 l0bl10 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b10c612 l0bl10 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b10c613 l0bl10 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b10c614 l0bl10 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b10c615 l0bl10 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b10c616 l0bl10 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b10c617 l0bl10 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b10c618 l0bl10 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b10c619 l0bl10 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b10c620 l0bl10 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b10c621 l0bl10 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b10c622 l0bl10 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b10c623 l0bl10 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b10c624 l0bl10 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b10c625 l0bl10 vdd x625 x625b CELLD r1=900e3 r0=10000e3
xl0b10c626 l0bl10 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b10c627 l0bl10 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b10c628 l0bl10 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b10c629 l0bl10 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b10c630 l0bl10 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b10c631 l0bl10 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b10c632 l0bl10 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b10c633 l0bl10 vdd x633 x633b CELLD r1=10000e3 r0=900e3
xl0b10c634 l0bl10 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b10c635 l0bl10 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b10c636 l0bl10 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b10c637 l0bl10 vdd x637 x637b CELLD r1=10000e3 r0=900e3
xl0b10c638 l0bl10 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b10c639 l0bl10 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b10c640 l0bl10 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b10c641 l0bl10 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b10c642 l0bl10 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b10c643 l0bl10 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b10c644 l0bl10 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b10c645 l0bl10 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b10c646 l0bl10 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b10c647 l0bl10 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b10c648 l0bl10 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b10c649 l0bl10 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b10c650 l0bl10 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b10c651 l0bl10 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b10c652 l0bl10 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b10c653 l0bl10 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b10c654 l0bl10 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b10c655 l0bl10 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b10c656 l0bl10 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b10c657 l0bl10 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b10c658 l0bl10 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b10c659 l0bl10 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b10c660 l0bl10 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b10c661 l0bl10 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b10c662 l0bl10 vdd x662 x662b CELLD r1=10000e3 r0=900e3
xl0b10c663 l0bl10 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b10c664 l0bl10 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b10c665 l0bl10 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b10c666 l0bl10 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b10c667 l0bl10 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b10c668 l0bl10 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b10c669 l0bl10 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b10c670 l0bl10 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b10c671 l0bl10 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b10c672 l0bl10 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b10c673 l0bl10 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b10c674 l0bl10 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b10c675 l0bl10 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b10c676 l0bl10 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b10c677 l0bl10 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b10c678 l0bl10 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b10c679 l0bl10 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b10c680 l0bl10 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b10c681 l0bl10 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b10c682 l0bl10 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b10c683 l0bl10 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b10c684 l0bl10 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b10c685 l0bl10 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b10c686 l0bl10 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b10c687 l0bl10 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b10c688 l0bl10 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b10c689 l0bl10 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b10c690 l0bl10 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b10c691 l0bl10 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b10c692 l0bl10 vdd x692 x692b CELLD r1=10000e3 r0=900e3
xl0b10c693 l0bl10 vdd x693 x693b CELLD r1=10000e3 r0=900e3
xl0b10c694 l0bl10 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b10c695 l0bl10 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b10c696 l0bl10 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b10c697 l0bl10 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b10c698 l0bl10 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b10c699 l0bl10 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b10c700 l0bl10 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b10c701 l0bl10 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b10c702 l0bl10 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b10c703 l0bl10 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b10c704 l0bl10 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b10c705 l0bl10 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b10c706 l0bl10 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b10c707 l0bl10 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b10c708 l0bl10 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b10c709 l0bl10 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b10c710 l0bl10 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b10c711 l0bl10 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b10c712 l0bl10 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b10c713 l0bl10 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b10c714 l0bl10 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b10c715 l0bl10 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b10c716 l0bl10 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b10c717 l0bl10 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b10c718 l0bl10 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b10c719 l0bl10 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b10c720 l0bl10 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b10c721 l0bl10 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b10c722 l0bl10 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b10c723 l0bl10 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b10c724 l0bl10 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b10c725 l0bl10 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b10c726 l0bl10 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b10c727 l0bl10 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b10c728 l0bl10 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b10c729 l0bl10 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b10c730 l0bl10 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b10c731 l0bl10 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b10c732 l0bl10 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b10c733 l0bl10 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b10c734 l0bl10 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b10c735 l0bl10 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b10c736 l0bl10 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b10c737 l0bl10 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b10c738 l0bl10 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b10c739 l0bl10 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b10c740 l0bl10 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b10c741 l0bl10 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b10c742 l0bl10 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b10c743 l0bl10 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b10c744 l0bl10 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b10c745 l0bl10 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b10c746 l0bl10 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b10c747 l0bl10 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b10c748 l0bl10 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b10c749 l0bl10 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b10c750 l0bl10 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b10c751 l0bl10 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b10c752 l0bl10 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b10c753 l0bl10 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b10c754 l0bl10 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b10c755 l0bl10 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b10c756 l0bl10 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b10c757 l0bl10 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b10c758 l0bl10 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b10c759 l0bl10 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b10c760 l0bl10 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b10c761 l0bl10 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b10c762 l0bl10 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b10c763 l0bl10 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b10c764 l0bl10 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b10c765 l0bl10 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b10c766 l0bl10 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b10c767 l0bl10 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b10c768 l0bl10 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b10c769 l0bl10 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b10c770 l0bl10 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b10c771 l0bl10 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b10c772 l0bl10 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b10c773 l0bl10 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b10c774 l0bl10 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b10c775 l0bl10 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b10c776 l0bl10 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b10c777 l0bl10 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b10c778 l0bl10 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b10c779 l0bl10 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b10c780 l0bl10 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b10c781 l0bl10 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b10c782 l0bl10 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b10c783 l0bl10 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b11c0 l0bl11 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b11c1 l0bl11 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b11c2 l0bl11 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b11c3 l0bl11 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b11c4 l0bl11 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b11c5 l0bl11 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b11c6 l0bl11 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b11c7 l0bl11 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b11c8 l0bl11 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b11c9 l0bl11 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b11c10 l0bl11 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b11c11 l0bl11 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b11c12 l0bl11 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b11c13 l0bl11 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b11c14 l0bl11 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b11c15 l0bl11 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b11c16 l0bl11 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b11c17 l0bl11 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b11c18 l0bl11 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b11c19 l0bl11 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b11c20 l0bl11 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b11c21 l0bl11 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b11c22 l0bl11 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b11c23 l0bl11 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b11c24 l0bl11 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b11c25 l0bl11 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b11c26 l0bl11 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b11c27 l0bl11 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b11c28 l0bl11 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b11c29 l0bl11 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b11c30 l0bl11 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b11c31 l0bl11 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b11c32 l0bl11 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b11c33 l0bl11 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b11c34 l0bl11 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b11c35 l0bl11 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b11c36 l0bl11 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b11c37 l0bl11 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b11c38 l0bl11 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b11c39 l0bl11 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b11c40 l0bl11 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b11c41 l0bl11 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b11c42 l0bl11 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b11c43 l0bl11 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b11c44 l0bl11 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b11c45 l0bl11 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b11c46 l0bl11 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b11c47 l0bl11 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b11c48 l0bl11 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b11c49 l0bl11 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b11c50 l0bl11 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b11c51 l0bl11 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b11c52 l0bl11 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b11c53 l0bl11 vdd x53 x53b CELLD r1=900e3 r0=10000e3
xl0b11c54 l0bl11 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b11c55 l0bl11 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b11c56 l0bl11 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b11c57 l0bl11 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b11c58 l0bl11 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b11c59 l0bl11 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b11c60 l0bl11 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b11c61 l0bl11 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b11c62 l0bl11 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b11c63 l0bl11 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b11c64 l0bl11 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b11c65 l0bl11 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b11c66 l0bl11 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b11c67 l0bl11 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b11c68 l0bl11 vdd x68 x68b CELLD r1=900e3 r0=10000e3
xl0b11c69 l0bl11 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b11c70 l0bl11 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b11c71 l0bl11 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b11c72 l0bl11 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b11c73 l0bl11 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b11c74 l0bl11 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b11c75 l0bl11 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b11c76 l0bl11 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b11c77 l0bl11 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b11c78 l0bl11 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b11c79 l0bl11 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b11c80 l0bl11 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b11c81 l0bl11 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b11c82 l0bl11 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b11c83 l0bl11 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b11c84 l0bl11 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b11c85 l0bl11 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b11c86 l0bl11 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b11c87 l0bl11 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b11c88 l0bl11 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b11c89 l0bl11 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b11c90 l0bl11 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b11c91 l0bl11 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b11c92 l0bl11 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b11c93 l0bl11 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b11c94 l0bl11 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b11c95 l0bl11 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b11c96 l0bl11 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b11c97 l0bl11 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b11c98 l0bl11 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b11c99 l0bl11 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b11c100 l0bl11 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b11c101 l0bl11 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b11c102 l0bl11 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b11c103 l0bl11 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b11c104 l0bl11 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b11c105 l0bl11 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b11c106 l0bl11 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b11c107 l0bl11 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b11c108 l0bl11 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b11c109 l0bl11 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b11c110 l0bl11 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b11c111 l0bl11 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b11c112 l0bl11 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b11c113 l0bl11 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b11c114 l0bl11 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b11c115 l0bl11 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b11c116 l0bl11 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b11c117 l0bl11 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b11c118 l0bl11 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b11c119 l0bl11 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b11c120 l0bl11 vdd x120 x120b CELLD r1=900e3 r0=10000e3
xl0b11c121 l0bl11 vdd x121 x121b CELLD r1=900e3 r0=10000e3
xl0b11c122 l0bl11 vdd x122 x122b CELLD r1=900e3 r0=10000e3
xl0b11c123 l0bl11 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b11c124 l0bl11 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b11c125 l0bl11 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b11c126 l0bl11 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b11c127 l0bl11 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b11c128 l0bl11 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b11c129 l0bl11 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b11c130 l0bl11 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b11c131 l0bl11 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b11c132 l0bl11 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b11c133 l0bl11 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b11c134 l0bl11 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b11c135 l0bl11 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b11c136 l0bl11 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b11c137 l0bl11 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b11c138 l0bl11 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b11c139 l0bl11 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b11c140 l0bl11 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b11c141 l0bl11 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b11c142 l0bl11 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b11c143 l0bl11 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b11c144 l0bl11 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b11c145 l0bl11 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b11c146 l0bl11 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b11c147 l0bl11 vdd x147 x147b CELLD r1=900e3 r0=10000e3
xl0b11c148 l0bl11 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b11c149 l0bl11 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b11c150 l0bl11 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b11c151 l0bl11 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b11c152 l0bl11 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b11c153 l0bl11 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b11c154 l0bl11 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b11c155 l0bl11 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b11c156 l0bl11 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b11c157 l0bl11 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b11c158 l0bl11 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b11c159 l0bl11 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b11c160 l0bl11 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b11c161 l0bl11 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b11c162 l0bl11 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b11c163 l0bl11 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b11c164 l0bl11 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b11c165 l0bl11 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b11c166 l0bl11 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b11c167 l0bl11 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b11c168 l0bl11 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b11c169 l0bl11 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b11c170 l0bl11 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b11c171 l0bl11 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b11c172 l0bl11 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b11c173 l0bl11 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b11c174 l0bl11 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b11c175 l0bl11 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b11c176 l0bl11 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b11c177 l0bl11 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b11c178 l0bl11 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b11c179 l0bl11 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b11c180 l0bl11 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b11c181 l0bl11 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b11c182 l0bl11 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b11c183 l0bl11 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b11c184 l0bl11 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b11c185 l0bl11 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b11c186 l0bl11 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b11c187 l0bl11 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b11c188 l0bl11 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b11c189 l0bl11 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b11c190 l0bl11 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b11c191 l0bl11 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b11c192 l0bl11 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b11c193 l0bl11 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b11c194 l0bl11 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b11c195 l0bl11 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b11c196 l0bl11 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b11c197 l0bl11 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b11c198 l0bl11 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b11c199 l0bl11 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b11c200 l0bl11 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b11c201 l0bl11 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b11c202 l0bl11 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b11c203 l0bl11 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b11c204 l0bl11 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b11c205 l0bl11 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b11c206 l0bl11 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b11c207 l0bl11 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b11c208 l0bl11 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b11c209 l0bl11 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b11c210 l0bl11 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b11c211 l0bl11 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b11c212 l0bl11 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b11c213 l0bl11 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b11c214 l0bl11 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b11c215 l0bl11 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b11c216 l0bl11 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b11c217 l0bl11 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b11c218 l0bl11 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b11c219 l0bl11 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b11c220 l0bl11 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b11c221 l0bl11 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b11c222 l0bl11 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b11c223 l0bl11 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b11c224 l0bl11 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b11c225 l0bl11 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b11c226 l0bl11 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b11c227 l0bl11 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b11c228 l0bl11 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b11c229 l0bl11 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b11c230 l0bl11 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b11c231 l0bl11 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b11c232 l0bl11 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b11c233 l0bl11 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b11c234 l0bl11 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b11c235 l0bl11 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b11c236 l0bl11 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b11c237 l0bl11 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b11c238 l0bl11 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b11c239 l0bl11 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b11c240 l0bl11 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b11c241 l0bl11 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b11c242 l0bl11 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b11c243 l0bl11 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b11c244 l0bl11 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b11c245 l0bl11 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b11c246 l0bl11 vdd x246 x246b CELLD r1=900e3 r0=10000e3
xl0b11c247 l0bl11 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b11c248 l0bl11 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b11c249 l0bl11 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b11c250 l0bl11 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b11c251 l0bl11 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b11c252 l0bl11 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b11c253 l0bl11 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b11c254 l0bl11 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b11c255 l0bl11 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b11c256 l0bl11 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b11c257 l0bl11 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b11c258 l0bl11 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b11c259 l0bl11 vdd x259 x259b CELLD r1=900e3 r0=10000e3
xl0b11c260 l0bl11 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b11c261 l0bl11 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b11c262 l0bl11 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b11c263 l0bl11 vdd x263 x263b CELLD r1=10000e3 r0=900e3
xl0b11c264 l0bl11 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b11c265 l0bl11 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b11c266 l0bl11 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b11c267 l0bl11 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b11c268 l0bl11 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b11c269 l0bl11 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b11c270 l0bl11 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b11c271 l0bl11 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b11c272 l0bl11 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b11c273 l0bl11 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b11c274 l0bl11 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b11c275 l0bl11 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b11c276 l0bl11 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b11c277 l0bl11 vdd x277 x277b CELLD r1=900e3 r0=10000e3
xl0b11c278 l0bl11 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b11c279 l0bl11 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b11c280 l0bl11 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b11c281 l0bl11 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b11c282 l0bl11 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b11c283 l0bl11 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b11c284 l0bl11 vdd x284 x284b CELLD r1=900e3 r0=10000e3
xl0b11c285 l0bl11 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b11c286 l0bl11 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b11c287 l0bl11 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b11c288 l0bl11 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b11c289 l0bl11 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b11c290 l0bl11 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b11c291 l0bl11 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b11c292 l0bl11 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b11c293 l0bl11 vdd x293 x293b CELLD r1=900e3 r0=10000e3
xl0b11c294 l0bl11 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b11c295 l0bl11 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b11c296 l0bl11 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b11c297 l0bl11 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b11c298 l0bl11 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b11c299 l0bl11 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b11c300 l0bl11 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b11c301 l0bl11 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b11c302 l0bl11 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b11c303 l0bl11 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b11c304 l0bl11 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b11c305 l0bl11 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b11c306 l0bl11 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b11c307 l0bl11 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b11c308 l0bl11 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b11c309 l0bl11 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b11c310 l0bl11 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b11c311 l0bl11 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b11c312 l0bl11 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b11c313 l0bl11 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b11c314 l0bl11 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b11c315 l0bl11 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b11c316 l0bl11 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b11c317 l0bl11 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b11c318 l0bl11 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b11c319 l0bl11 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b11c320 l0bl11 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b11c321 l0bl11 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b11c322 l0bl11 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b11c323 l0bl11 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b11c324 l0bl11 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b11c325 l0bl11 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b11c326 l0bl11 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b11c327 l0bl11 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b11c328 l0bl11 vdd x328 x328b CELLD r1=900e3 r0=10000e3
xl0b11c329 l0bl11 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b11c330 l0bl11 vdd x330 x330b CELLD r1=900e3 r0=10000e3
xl0b11c331 l0bl11 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b11c332 l0bl11 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b11c333 l0bl11 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b11c334 l0bl11 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b11c335 l0bl11 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b11c336 l0bl11 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b11c337 l0bl11 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b11c338 l0bl11 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b11c339 l0bl11 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b11c340 l0bl11 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b11c341 l0bl11 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b11c342 l0bl11 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b11c343 l0bl11 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b11c344 l0bl11 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b11c345 l0bl11 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b11c346 l0bl11 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b11c347 l0bl11 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b11c348 l0bl11 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b11c349 l0bl11 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b11c350 l0bl11 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b11c351 l0bl11 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b11c352 l0bl11 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b11c353 l0bl11 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b11c354 l0bl11 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b11c355 l0bl11 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b11c356 l0bl11 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b11c357 l0bl11 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b11c358 l0bl11 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b11c359 l0bl11 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b11c360 l0bl11 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b11c361 l0bl11 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b11c362 l0bl11 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b11c363 l0bl11 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b11c364 l0bl11 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b11c365 l0bl11 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b11c366 l0bl11 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b11c367 l0bl11 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b11c368 l0bl11 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b11c369 l0bl11 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b11c370 l0bl11 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b11c371 l0bl11 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b11c372 l0bl11 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b11c373 l0bl11 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b11c374 l0bl11 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b11c375 l0bl11 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b11c376 l0bl11 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b11c377 l0bl11 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b11c378 l0bl11 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b11c379 l0bl11 vdd x379 x379b CELLD r1=10000e3 r0=900e3
xl0b11c380 l0bl11 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b11c381 l0bl11 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b11c382 l0bl11 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b11c383 l0bl11 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b11c384 l0bl11 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b11c385 l0bl11 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b11c386 l0bl11 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b11c387 l0bl11 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b11c388 l0bl11 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b11c389 l0bl11 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b11c390 l0bl11 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b11c391 l0bl11 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b11c392 l0bl11 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b11c393 l0bl11 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b11c394 l0bl11 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b11c395 l0bl11 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b11c396 l0bl11 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b11c397 l0bl11 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b11c398 l0bl11 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b11c399 l0bl11 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b11c400 l0bl11 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b11c401 l0bl11 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b11c402 l0bl11 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b11c403 l0bl11 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b11c404 l0bl11 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b11c405 l0bl11 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b11c406 l0bl11 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b11c407 l0bl11 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b11c408 l0bl11 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b11c409 l0bl11 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b11c410 l0bl11 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b11c411 l0bl11 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b11c412 l0bl11 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b11c413 l0bl11 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b11c414 l0bl11 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b11c415 l0bl11 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b11c416 l0bl11 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b11c417 l0bl11 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b11c418 l0bl11 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b11c419 l0bl11 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b11c420 l0bl11 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b11c421 l0bl11 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b11c422 l0bl11 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b11c423 l0bl11 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b11c424 l0bl11 vdd x424 x424b CELLD r1=900e3 r0=10000e3
xl0b11c425 l0bl11 vdd x425 x425b CELLD r1=900e3 r0=10000e3
xl0b11c426 l0bl11 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b11c427 l0bl11 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b11c428 l0bl11 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b11c429 l0bl11 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b11c430 l0bl11 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b11c431 l0bl11 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b11c432 l0bl11 vdd x432 x432b CELLD r1=10000e3 r0=900e3
xl0b11c433 l0bl11 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b11c434 l0bl11 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b11c435 l0bl11 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b11c436 l0bl11 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b11c437 l0bl11 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b11c438 l0bl11 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b11c439 l0bl11 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b11c440 l0bl11 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b11c441 l0bl11 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b11c442 l0bl11 vdd x442 x442b CELLD r1=900e3 r0=10000e3
xl0b11c443 l0bl11 vdd x443 x443b CELLD r1=900e3 r0=10000e3
xl0b11c444 l0bl11 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b11c445 l0bl11 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b11c446 l0bl11 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b11c447 l0bl11 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b11c448 l0bl11 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b11c449 l0bl11 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b11c450 l0bl11 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b11c451 l0bl11 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b11c452 l0bl11 vdd x452 x452b CELLD r1=900e3 r0=10000e3
xl0b11c453 l0bl11 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b11c454 l0bl11 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b11c455 l0bl11 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b11c456 l0bl11 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b11c457 l0bl11 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b11c458 l0bl11 vdd x458 x458b CELLD r1=10000e3 r0=900e3
xl0b11c459 l0bl11 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b11c460 l0bl11 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b11c461 l0bl11 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b11c462 l0bl11 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b11c463 l0bl11 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b11c464 l0bl11 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b11c465 l0bl11 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b11c466 l0bl11 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b11c467 l0bl11 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b11c468 l0bl11 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b11c469 l0bl11 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b11c470 l0bl11 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b11c471 l0bl11 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b11c472 l0bl11 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b11c473 l0bl11 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b11c474 l0bl11 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b11c475 l0bl11 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b11c476 l0bl11 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b11c477 l0bl11 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b11c478 l0bl11 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b11c479 l0bl11 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b11c480 l0bl11 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b11c481 l0bl11 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b11c482 l0bl11 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b11c483 l0bl11 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b11c484 l0bl11 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b11c485 l0bl11 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b11c486 l0bl11 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b11c487 l0bl11 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b11c488 l0bl11 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b11c489 l0bl11 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b11c490 l0bl11 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b11c491 l0bl11 vdd x491 x491b CELLD r1=10000e3 r0=900e3
xl0b11c492 l0bl11 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b11c493 l0bl11 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b11c494 l0bl11 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b11c495 l0bl11 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b11c496 l0bl11 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b11c497 l0bl11 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b11c498 l0bl11 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b11c499 l0bl11 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b11c500 l0bl11 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b11c501 l0bl11 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b11c502 l0bl11 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b11c503 l0bl11 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b11c504 l0bl11 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b11c505 l0bl11 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b11c506 l0bl11 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b11c507 l0bl11 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b11c508 l0bl11 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b11c509 l0bl11 vdd x509 x509b CELLD r1=900e3 r0=10000e3
xl0b11c510 l0bl11 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b11c511 l0bl11 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b11c512 l0bl11 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b11c513 l0bl11 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b11c514 l0bl11 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b11c515 l0bl11 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b11c516 l0bl11 vdd x516 x516b CELLD r1=10000e3 r0=900e3
xl0b11c517 l0bl11 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b11c518 l0bl11 vdd x518 x518b CELLD r1=10000e3 r0=900e3
xl0b11c519 l0bl11 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b11c520 l0bl11 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b11c521 l0bl11 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b11c522 l0bl11 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b11c523 l0bl11 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b11c524 l0bl11 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b11c525 l0bl11 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b11c526 l0bl11 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b11c527 l0bl11 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b11c528 l0bl11 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b11c529 l0bl11 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b11c530 l0bl11 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b11c531 l0bl11 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b11c532 l0bl11 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b11c533 l0bl11 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b11c534 l0bl11 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b11c535 l0bl11 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b11c536 l0bl11 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b11c537 l0bl11 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b11c538 l0bl11 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b11c539 l0bl11 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b11c540 l0bl11 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b11c541 l0bl11 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b11c542 l0bl11 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b11c543 l0bl11 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b11c544 l0bl11 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b11c545 l0bl11 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b11c546 l0bl11 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b11c547 l0bl11 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b11c548 l0bl11 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b11c549 l0bl11 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b11c550 l0bl11 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b11c551 l0bl11 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b11c552 l0bl11 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b11c553 l0bl11 vdd x553 x553b CELLD r1=900e3 r0=10000e3
xl0b11c554 l0bl11 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b11c555 l0bl11 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b11c556 l0bl11 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b11c557 l0bl11 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b11c558 l0bl11 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b11c559 l0bl11 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b11c560 l0bl11 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b11c561 l0bl11 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b11c562 l0bl11 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b11c563 l0bl11 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b11c564 l0bl11 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b11c565 l0bl11 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b11c566 l0bl11 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b11c567 l0bl11 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b11c568 l0bl11 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b11c569 l0bl11 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b11c570 l0bl11 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b11c571 l0bl11 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b11c572 l0bl11 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b11c573 l0bl11 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b11c574 l0bl11 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b11c575 l0bl11 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b11c576 l0bl11 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b11c577 l0bl11 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b11c578 l0bl11 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b11c579 l0bl11 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b11c580 l0bl11 vdd x580 x580b CELLD r1=900e3 r0=10000e3
xl0b11c581 l0bl11 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b11c582 l0bl11 vdd x582 x582b CELLD r1=900e3 r0=10000e3
xl0b11c583 l0bl11 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b11c584 l0bl11 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b11c585 l0bl11 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b11c586 l0bl11 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b11c587 l0bl11 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b11c588 l0bl11 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b11c589 l0bl11 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b11c590 l0bl11 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b11c591 l0bl11 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b11c592 l0bl11 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b11c593 l0bl11 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b11c594 l0bl11 vdd x594 x594b CELLD r1=900e3 r0=10000e3
xl0b11c595 l0bl11 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b11c596 l0bl11 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b11c597 l0bl11 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b11c598 l0bl11 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b11c599 l0bl11 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b11c600 l0bl11 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b11c601 l0bl11 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b11c602 l0bl11 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b11c603 l0bl11 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b11c604 l0bl11 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b11c605 l0bl11 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b11c606 l0bl11 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b11c607 l0bl11 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b11c608 l0bl11 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b11c609 l0bl11 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b11c610 l0bl11 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b11c611 l0bl11 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b11c612 l0bl11 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b11c613 l0bl11 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b11c614 l0bl11 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b11c615 l0bl11 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b11c616 l0bl11 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b11c617 l0bl11 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b11c618 l0bl11 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b11c619 l0bl11 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b11c620 l0bl11 vdd x620 x620b CELLD r1=900e3 r0=10000e3
xl0b11c621 l0bl11 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b11c622 l0bl11 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b11c623 l0bl11 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b11c624 l0bl11 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b11c625 l0bl11 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b11c626 l0bl11 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b11c627 l0bl11 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b11c628 l0bl11 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b11c629 l0bl11 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b11c630 l0bl11 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b11c631 l0bl11 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b11c632 l0bl11 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b11c633 l0bl11 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b11c634 l0bl11 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b11c635 l0bl11 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b11c636 l0bl11 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b11c637 l0bl11 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b11c638 l0bl11 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b11c639 l0bl11 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b11c640 l0bl11 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b11c641 l0bl11 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b11c642 l0bl11 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b11c643 l0bl11 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b11c644 l0bl11 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b11c645 l0bl11 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b11c646 l0bl11 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b11c647 l0bl11 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b11c648 l0bl11 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b11c649 l0bl11 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b11c650 l0bl11 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b11c651 l0bl11 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b11c652 l0bl11 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b11c653 l0bl11 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b11c654 l0bl11 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b11c655 l0bl11 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b11c656 l0bl11 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b11c657 l0bl11 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b11c658 l0bl11 vdd x658 x658b CELLD r1=900e3 r0=10000e3
xl0b11c659 l0bl11 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b11c660 l0bl11 vdd x660 x660b CELLD r1=900e3 r0=10000e3
xl0b11c661 l0bl11 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b11c662 l0bl11 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b11c663 l0bl11 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b11c664 l0bl11 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b11c665 l0bl11 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b11c666 l0bl11 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b11c667 l0bl11 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b11c668 l0bl11 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b11c669 l0bl11 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b11c670 l0bl11 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b11c671 l0bl11 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b11c672 l0bl11 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b11c673 l0bl11 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b11c674 l0bl11 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b11c675 l0bl11 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b11c676 l0bl11 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b11c677 l0bl11 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b11c678 l0bl11 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b11c679 l0bl11 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b11c680 l0bl11 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b11c681 l0bl11 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b11c682 l0bl11 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b11c683 l0bl11 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b11c684 l0bl11 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b11c685 l0bl11 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b11c686 l0bl11 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b11c687 l0bl11 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b11c688 l0bl11 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b11c689 l0bl11 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b11c690 l0bl11 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b11c691 l0bl11 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b11c692 l0bl11 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b11c693 l0bl11 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b11c694 l0bl11 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b11c695 l0bl11 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b11c696 l0bl11 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b11c697 l0bl11 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b11c698 l0bl11 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b11c699 l0bl11 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b11c700 l0bl11 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b11c701 l0bl11 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b11c702 l0bl11 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b11c703 l0bl11 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b11c704 l0bl11 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b11c705 l0bl11 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b11c706 l0bl11 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b11c707 l0bl11 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b11c708 l0bl11 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b11c709 l0bl11 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b11c710 l0bl11 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b11c711 l0bl11 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b11c712 l0bl11 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b11c713 l0bl11 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b11c714 l0bl11 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b11c715 l0bl11 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b11c716 l0bl11 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b11c717 l0bl11 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b11c718 l0bl11 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b11c719 l0bl11 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b11c720 l0bl11 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b11c721 l0bl11 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b11c722 l0bl11 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b11c723 l0bl11 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b11c724 l0bl11 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b11c725 l0bl11 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b11c726 l0bl11 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b11c727 l0bl11 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b11c728 l0bl11 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b11c729 l0bl11 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b11c730 l0bl11 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b11c731 l0bl11 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b11c732 l0bl11 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b11c733 l0bl11 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b11c734 l0bl11 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b11c735 l0bl11 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b11c736 l0bl11 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b11c737 l0bl11 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b11c738 l0bl11 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b11c739 l0bl11 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b11c740 l0bl11 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b11c741 l0bl11 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b11c742 l0bl11 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b11c743 l0bl11 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b11c744 l0bl11 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b11c745 l0bl11 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b11c746 l0bl11 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b11c747 l0bl11 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b11c748 l0bl11 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b11c749 l0bl11 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b11c750 l0bl11 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b11c751 l0bl11 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b11c752 l0bl11 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b11c753 l0bl11 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b11c754 l0bl11 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b11c755 l0bl11 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b11c756 l0bl11 vdd x756 x756b CELLD r1=900e3 r0=10000e3
xl0b11c757 l0bl11 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b11c758 l0bl11 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b11c759 l0bl11 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b11c760 l0bl11 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b11c761 l0bl11 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b11c762 l0bl11 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b11c763 l0bl11 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b11c764 l0bl11 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b11c765 l0bl11 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b11c766 l0bl11 vdd x766 x766b CELLD r1=900e3 r0=10000e3
xl0b11c767 l0bl11 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b11c768 l0bl11 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b11c769 l0bl11 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b11c770 l0bl11 vdd x770 x770b CELLD r1=900e3 r0=10000e3
xl0b11c771 l0bl11 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b11c772 l0bl11 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b11c773 l0bl11 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b11c774 l0bl11 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b11c775 l0bl11 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b11c776 l0bl11 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b11c777 l0bl11 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b11c778 l0bl11 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b11c779 l0bl11 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b11c780 l0bl11 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b11c781 l0bl11 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b11c782 l0bl11 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b11c783 l0bl11 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b12c0 l0bl12 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b12c1 l0bl12 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b12c2 l0bl12 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b12c3 l0bl12 vdd x3 x3b CELLD r1=10000e3 r0=900e3
xl0b12c4 l0bl12 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b12c5 l0bl12 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b12c6 l0bl12 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b12c7 l0bl12 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b12c8 l0bl12 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b12c9 l0bl12 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b12c10 l0bl12 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b12c11 l0bl12 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b12c12 l0bl12 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b12c13 l0bl12 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b12c14 l0bl12 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b12c15 l0bl12 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b12c16 l0bl12 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b12c17 l0bl12 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b12c18 l0bl12 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b12c19 l0bl12 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b12c20 l0bl12 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b12c21 l0bl12 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b12c22 l0bl12 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b12c23 l0bl12 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b12c24 l0bl12 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b12c25 l0bl12 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b12c26 l0bl12 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b12c27 l0bl12 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b12c28 l0bl12 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b12c29 l0bl12 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b12c30 l0bl12 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b12c31 l0bl12 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b12c32 l0bl12 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b12c33 l0bl12 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b12c34 l0bl12 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b12c35 l0bl12 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b12c36 l0bl12 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b12c37 l0bl12 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b12c38 l0bl12 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b12c39 l0bl12 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b12c40 l0bl12 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b12c41 l0bl12 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b12c42 l0bl12 vdd x42 x42b CELLD r1=10000e3 r0=900e3
xl0b12c43 l0bl12 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b12c44 l0bl12 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b12c45 l0bl12 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b12c46 l0bl12 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b12c47 l0bl12 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b12c48 l0bl12 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b12c49 l0bl12 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b12c50 l0bl12 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b12c51 l0bl12 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b12c52 l0bl12 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b12c53 l0bl12 vdd x53 x53b CELLD r1=900e3 r0=10000e3
xl0b12c54 l0bl12 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b12c55 l0bl12 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b12c56 l0bl12 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b12c57 l0bl12 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b12c58 l0bl12 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b12c59 l0bl12 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b12c60 l0bl12 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b12c61 l0bl12 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b12c62 l0bl12 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b12c63 l0bl12 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b12c64 l0bl12 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b12c65 l0bl12 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b12c66 l0bl12 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b12c67 l0bl12 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b12c68 l0bl12 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b12c69 l0bl12 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b12c70 l0bl12 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b12c71 l0bl12 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b12c72 l0bl12 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b12c73 l0bl12 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b12c74 l0bl12 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b12c75 l0bl12 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b12c76 l0bl12 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b12c77 l0bl12 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b12c78 l0bl12 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b12c79 l0bl12 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b12c80 l0bl12 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b12c81 l0bl12 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b12c82 l0bl12 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b12c83 l0bl12 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b12c84 l0bl12 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b12c85 l0bl12 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b12c86 l0bl12 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b12c87 l0bl12 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b12c88 l0bl12 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b12c89 l0bl12 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b12c90 l0bl12 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b12c91 l0bl12 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b12c92 l0bl12 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b12c93 l0bl12 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b12c94 l0bl12 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b12c95 l0bl12 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b12c96 l0bl12 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b12c97 l0bl12 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b12c98 l0bl12 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b12c99 l0bl12 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b12c100 l0bl12 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b12c101 l0bl12 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b12c102 l0bl12 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b12c103 l0bl12 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b12c104 l0bl12 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b12c105 l0bl12 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b12c106 l0bl12 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b12c107 l0bl12 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b12c108 l0bl12 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b12c109 l0bl12 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b12c110 l0bl12 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b12c111 l0bl12 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b12c112 l0bl12 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b12c113 l0bl12 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b12c114 l0bl12 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b12c115 l0bl12 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b12c116 l0bl12 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b12c117 l0bl12 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b12c118 l0bl12 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b12c119 l0bl12 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b12c120 l0bl12 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b12c121 l0bl12 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b12c122 l0bl12 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b12c123 l0bl12 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b12c124 l0bl12 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b12c125 l0bl12 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b12c126 l0bl12 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b12c127 l0bl12 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b12c128 l0bl12 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b12c129 l0bl12 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b12c130 l0bl12 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b12c131 l0bl12 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b12c132 l0bl12 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b12c133 l0bl12 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b12c134 l0bl12 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b12c135 l0bl12 vdd x135 x135b CELLD r1=900e3 r0=10000e3
xl0b12c136 l0bl12 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b12c137 l0bl12 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b12c138 l0bl12 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b12c139 l0bl12 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b12c140 l0bl12 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b12c141 l0bl12 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b12c142 l0bl12 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b12c143 l0bl12 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b12c144 l0bl12 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b12c145 l0bl12 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b12c146 l0bl12 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b12c147 l0bl12 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b12c148 l0bl12 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b12c149 l0bl12 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b12c150 l0bl12 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b12c151 l0bl12 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b12c152 l0bl12 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b12c153 l0bl12 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b12c154 l0bl12 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b12c155 l0bl12 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b12c156 l0bl12 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b12c157 l0bl12 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b12c158 l0bl12 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b12c159 l0bl12 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b12c160 l0bl12 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b12c161 l0bl12 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b12c162 l0bl12 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b12c163 l0bl12 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b12c164 l0bl12 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b12c165 l0bl12 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b12c166 l0bl12 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b12c167 l0bl12 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b12c168 l0bl12 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b12c169 l0bl12 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b12c170 l0bl12 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b12c171 l0bl12 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b12c172 l0bl12 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b12c173 l0bl12 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b12c174 l0bl12 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b12c175 l0bl12 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b12c176 l0bl12 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b12c177 l0bl12 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b12c178 l0bl12 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b12c179 l0bl12 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b12c180 l0bl12 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b12c181 l0bl12 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b12c182 l0bl12 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b12c183 l0bl12 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b12c184 l0bl12 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b12c185 l0bl12 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b12c186 l0bl12 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b12c187 l0bl12 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b12c188 l0bl12 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b12c189 l0bl12 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b12c190 l0bl12 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b12c191 l0bl12 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b12c192 l0bl12 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b12c193 l0bl12 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b12c194 l0bl12 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b12c195 l0bl12 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b12c196 l0bl12 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b12c197 l0bl12 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b12c198 l0bl12 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b12c199 l0bl12 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b12c200 l0bl12 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b12c201 l0bl12 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b12c202 l0bl12 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b12c203 l0bl12 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b12c204 l0bl12 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b12c205 l0bl12 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b12c206 l0bl12 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b12c207 l0bl12 vdd x207 x207b CELLD r1=900e3 r0=10000e3
xl0b12c208 l0bl12 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b12c209 l0bl12 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b12c210 l0bl12 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b12c211 l0bl12 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b12c212 l0bl12 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b12c213 l0bl12 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b12c214 l0bl12 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b12c215 l0bl12 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b12c216 l0bl12 vdd x216 x216b CELLD r1=900e3 r0=10000e3
xl0b12c217 l0bl12 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b12c218 l0bl12 vdd x218 x218b CELLD r1=900e3 r0=10000e3
xl0b12c219 l0bl12 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b12c220 l0bl12 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b12c221 l0bl12 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b12c222 l0bl12 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b12c223 l0bl12 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b12c224 l0bl12 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b12c225 l0bl12 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b12c226 l0bl12 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b12c227 l0bl12 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b12c228 l0bl12 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b12c229 l0bl12 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b12c230 l0bl12 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b12c231 l0bl12 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b12c232 l0bl12 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b12c233 l0bl12 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b12c234 l0bl12 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b12c235 l0bl12 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b12c236 l0bl12 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b12c237 l0bl12 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b12c238 l0bl12 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b12c239 l0bl12 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b12c240 l0bl12 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b12c241 l0bl12 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b12c242 l0bl12 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b12c243 l0bl12 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b12c244 l0bl12 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b12c245 l0bl12 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b12c246 l0bl12 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b12c247 l0bl12 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b12c248 l0bl12 vdd x248 x248b CELLD r1=900e3 r0=10000e3
xl0b12c249 l0bl12 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b12c250 l0bl12 vdd x250 x250b CELLD r1=900e3 r0=10000e3
xl0b12c251 l0bl12 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b12c252 l0bl12 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b12c253 l0bl12 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b12c254 l0bl12 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b12c255 l0bl12 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b12c256 l0bl12 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b12c257 l0bl12 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b12c258 l0bl12 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b12c259 l0bl12 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b12c260 l0bl12 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b12c261 l0bl12 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b12c262 l0bl12 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b12c263 l0bl12 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b12c264 l0bl12 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b12c265 l0bl12 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b12c266 l0bl12 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b12c267 l0bl12 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b12c268 l0bl12 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b12c269 l0bl12 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b12c270 l0bl12 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b12c271 l0bl12 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b12c272 l0bl12 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b12c273 l0bl12 vdd x273 x273b CELLD r1=900e3 r0=10000e3
xl0b12c274 l0bl12 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b12c275 l0bl12 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b12c276 l0bl12 vdd x276 x276b CELLD r1=900e3 r0=10000e3
xl0b12c277 l0bl12 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b12c278 l0bl12 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b12c279 l0bl12 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b12c280 l0bl12 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b12c281 l0bl12 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b12c282 l0bl12 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b12c283 l0bl12 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b12c284 l0bl12 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b12c285 l0bl12 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b12c286 l0bl12 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b12c287 l0bl12 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b12c288 l0bl12 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b12c289 l0bl12 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b12c290 l0bl12 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b12c291 l0bl12 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b12c292 l0bl12 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b12c293 l0bl12 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b12c294 l0bl12 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b12c295 l0bl12 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b12c296 l0bl12 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b12c297 l0bl12 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b12c298 l0bl12 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b12c299 l0bl12 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b12c300 l0bl12 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b12c301 l0bl12 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b12c302 l0bl12 vdd x302 x302b CELLD r1=900e3 r0=10000e3
xl0b12c303 l0bl12 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b12c304 l0bl12 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b12c305 l0bl12 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b12c306 l0bl12 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b12c307 l0bl12 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b12c308 l0bl12 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b12c309 l0bl12 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b12c310 l0bl12 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b12c311 l0bl12 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b12c312 l0bl12 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b12c313 l0bl12 vdd x313 x313b CELLD r1=900e3 r0=10000e3
xl0b12c314 l0bl12 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b12c315 l0bl12 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b12c316 l0bl12 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b12c317 l0bl12 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b12c318 l0bl12 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b12c319 l0bl12 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b12c320 l0bl12 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b12c321 l0bl12 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b12c322 l0bl12 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b12c323 l0bl12 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b12c324 l0bl12 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b12c325 l0bl12 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b12c326 l0bl12 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b12c327 l0bl12 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b12c328 l0bl12 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b12c329 l0bl12 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b12c330 l0bl12 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b12c331 l0bl12 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b12c332 l0bl12 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b12c333 l0bl12 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b12c334 l0bl12 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b12c335 l0bl12 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b12c336 l0bl12 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b12c337 l0bl12 vdd x337 x337b CELLD r1=10000e3 r0=900e3
xl0b12c338 l0bl12 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b12c339 l0bl12 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b12c340 l0bl12 vdd x340 x340b CELLD r1=900e3 r0=10000e3
xl0b12c341 l0bl12 vdd x341 x341b CELLD r1=900e3 r0=10000e3
xl0b12c342 l0bl12 vdd x342 x342b CELLD r1=900e3 r0=10000e3
xl0b12c343 l0bl12 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b12c344 l0bl12 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b12c345 l0bl12 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b12c346 l0bl12 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b12c347 l0bl12 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b12c348 l0bl12 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b12c349 l0bl12 vdd x349 x349b CELLD r1=10000e3 r0=900e3
xl0b12c350 l0bl12 vdd x350 x350b CELLD r1=10000e3 r0=900e3
xl0b12c351 l0bl12 vdd x351 x351b CELLD r1=10000e3 r0=900e3
xl0b12c352 l0bl12 vdd x352 x352b CELLD r1=10000e3 r0=900e3
xl0b12c353 l0bl12 vdd x353 x353b CELLD r1=10000e3 r0=900e3
xl0b12c354 l0bl12 vdd x354 x354b CELLD r1=10000e3 r0=900e3
xl0b12c355 l0bl12 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b12c356 l0bl12 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b12c357 l0bl12 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b12c358 l0bl12 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b12c359 l0bl12 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b12c360 l0bl12 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b12c361 l0bl12 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b12c362 l0bl12 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b12c363 l0bl12 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b12c364 l0bl12 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b12c365 l0bl12 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b12c366 l0bl12 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b12c367 l0bl12 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b12c368 l0bl12 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b12c369 l0bl12 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b12c370 l0bl12 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b12c371 l0bl12 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b12c372 l0bl12 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b12c373 l0bl12 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b12c374 l0bl12 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b12c375 l0bl12 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b12c376 l0bl12 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b12c377 l0bl12 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b12c378 l0bl12 vdd x378 x378b CELLD r1=10000e3 r0=900e3
xl0b12c379 l0bl12 vdd x379 x379b CELLD r1=10000e3 r0=900e3
xl0b12c380 l0bl12 vdd x380 x380b CELLD r1=10000e3 r0=900e3
xl0b12c381 l0bl12 vdd x381 x381b CELLD r1=10000e3 r0=900e3
xl0b12c382 l0bl12 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b12c383 l0bl12 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b12c384 l0bl12 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b12c385 l0bl12 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b12c386 l0bl12 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b12c387 l0bl12 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b12c388 l0bl12 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b12c389 l0bl12 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b12c390 l0bl12 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b12c391 l0bl12 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b12c392 l0bl12 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b12c393 l0bl12 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b12c394 l0bl12 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b12c395 l0bl12 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b12c396 l0bl12 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b12c397 l0bl12 vdd x397 x397b CELLD r1=900e3 r0=10000e3
xl0b12c398 l0bl12 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b12c399 l0bl12 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b12c400 l0bl12 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b12c401 l0bl12 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b12c402 l0bl12 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b12c403 l0bl12 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b12c404 l0bl12 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b12c405 l0bl12 vdd x405 x405b CELLD r1=10000e3 r0=900e3
xl0b12c406 l0bl12 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b12c407 l0bl12 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b12c408 l0bl12 vdd x408 x408b CELLD r1=10000e3 r0=900e3
xl0b12c409 l0bl12 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b12c410 l0bl12 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b12c411 l0bl12 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b12c412 l0bl12 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b12c413 l0bl12 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b12c414 l0bl12 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b12c415 l0bl12 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b12c416 l0bl12 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b12c417 l0bl12 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b12c418 l0bl12 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b12c419 l0bl12 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b12c420 l0bl12 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b12c421 l0bl12 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b12c422 l0bl12 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b12c423 l0bl12 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b12c424 l0bl12 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b12c425 l0bl12 vdd x425 x425b CELLD r1=900e3 r0=10000e3
xl0b12c426 l0bl12 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b12c427 l0bl12 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b12c428 l0bl12 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b12c429 l0bl12 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b12c430 l0bl12 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b12c431 l0bl12 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b12c432 l0bl12 vdd x432 x432b CELLD r1=10000e3 r0=900e3
xl0b12c433 l0bl12 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b12c434 l0bl12 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b12c435 l0bl12 vdd x435 x435b CELLD r1=10000e3 r0=900e3
xl0b12c436 l0bl12 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b12c437 l0bl12 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b12c438 l0bl12 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b12c439 l0bl12 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b12c440 l0bl12 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b12c441 l0bl12 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b12c442 l0bl12 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b12c443 l0bl12 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b12c444 l0bl12 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b12c445 l0bl12 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b12c446 l0bl12 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b12c447 l0bl12 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b12c448 l0bl12 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b12c449 l0bl12 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b12c450 l0bl12 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b12c451 l0bl12 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b12c452 l0bl12 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b12c453 l0bl12 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b12c454 l0bl12 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b12c455 l0bl12 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b12c456 l0bl12 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b12c457 l0bl12 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b12c458 l0bl12 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b12c459 l0bl12 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b12c460 l0bl12 vdd x460 x460b CELLD r1=10000e3 r0=900e3
xl0b12c461 l0bl12 vdd x461 x461b CELLD r1=10000e3 r0=900e3
xl0b12c462 l0bl12 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b12c463 l0bl12 vdd x463 x463b CELLD r1=10000e3 r0=900e3
xl0b12c464 l0bl12 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b12c465 l0bl12 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b12c466 l0bl12 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b12c467 l0bl12 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b12c468 l0bl12 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b12c469 l0bl12 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b12c470 l0bl12 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b12c471 l0bl12 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b12c472 l0bl12 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b12c473 l0bl12 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b12c474 l0bl12 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b12c475 l0bl12 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b12c476 l0bl12 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b12c477 l0bl12 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b12c478 l0bl12 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b12c479 l0bl12 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b12c480 l0bl12 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b12c481 l0bl12 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b12c482 l0bl12 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b12c483 l0bl12 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b12c484 l0bl12 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b12c485 l0bl12 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b12c486 l0bl12 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b12c487 l0bl12 vdd x487 x487b CELLD r1=10000e3 r0=900e3
xl0b12c488 l0bl12 vdd x488 x488b CELLD r1=10000e3 r0=900e3
xl0b12c489 l0bl12 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b12c490 l0bl12 vdd x490 x490b CELLD r1=10000e3 r0=900e3
xl0b12c491 l0bl12 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b12c492 l0bl12 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b12c493 l0bl12 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b12c494 l0bl12 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b12c495 l0bl12 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b12c496 l0bl12 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b12c497 l0bl12 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b12c498 l0bl12 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b12c499 l0bl12 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b12c500 l0bl12 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b12c501 l0bl12 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b12c502 l0bl12 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b12c503 l0bl12 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b12c504 l0bl12 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b12c505 l0bl12 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b12c506 l0bl12 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b12c507 l0bl12 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b12c508 l0bl12 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b12c509 l0bl12 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b12c510 l0bl12 vdd x510 x510b CELLD r1=900e3 r0=10000e3
xl0b12c511 l0bl12 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b12c512 l0bl12 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b12c513 l0bl12 vdd x513 x513b CELLD r1=10000e3 r0=900e3
xl0b12c514 l0bl12 vdd x514 x514b CELLD r1=10000e3 r0=900e3
xl0b12c515 l0bl12 vdd x515 x515b CELLD r1=10000e3 r0=900e3
xl0b12c516 l0bl12 vdd x516 x516b CELLD r1=10000e3 r0=900e3
xl0b12c517 l0bl12 vdd x517 x517b CELLD r1=10000e3 r0=900e3
xl0b12c518 l0bl12 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b12c519 l0bl12 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b12c520 l0bl12 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b12c521 l0bl12 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b12c522 l0bl12 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b12c523 l0bl12 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b12c524 l0bl12 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b12c525 l0bl12 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b12c526 l0bl12 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b12c527 l0bl12 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b12c528 l0bl12 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b12c529 l0bl12 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b12c530 l0bl12 vdd x530 x530b CELLD r1=10000e3 r0=900e3
xl0b12c531 l0bl12 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b12c532 l0bl12 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b12c533 l0bl12 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b12c534 l0bl12 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b12c535 l0bl12 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b12c536 l0bl12 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b12c537 l0bl12 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b12c538 l0bl12 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b12c539 l0bl12 vdd x539 x539b CELLD r1=900e3 r0=10000e3
xl0b12c540 l0bl12 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b12c541 l0bl12 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b12c542 l0bl12 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b12c543 l0bl12 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b12c544 l0bl12 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b12c545 l0bl12 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b12c546 l0bl12 vdd x546 x546b CELLD r1=10000e3 r0=900e3
xl0b12c547 l0bl12 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b12c548 l0bl12 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b12c549 l0bl12 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b12c550 l0bl12 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b12c551 l0bl12 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b12c552 l0bl12 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b12c553 l0bl12 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b12c554 l0bl12 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b12c555 l0bl12 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b12c556 l0bl12 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b12c557 l0bl12 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b12c558 l0bl12 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b12c559 l0bl12 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b12c560 l0bl12 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b12c561 l0bl12 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b12c562 l0bl12 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b12c563 l0bl12 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b12c564 l0bl12 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b12c565 l0bl12 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b12c566 l0bl12 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b12c567 l0bl12 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b12c568 l0bl12 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b12c569 l0bl12 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b12c570 l0bl12 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b12c571 l0bl12 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b12c572 l0bl12 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b12c573 l0bl12 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b12c574 l0bl12 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b12c575 l0bl12 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b12c576 l0bl12 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b12c577 l0bl12 vdd x577 x577b CELLD r1=10000e3 r0=900e3
xl0b12c578 l0bl12 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b12c579 l0bl12 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b12c580 l0bl12 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b12c581 l0bl12 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b12c582 l0bl12 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b12c583 l0bl12 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b12c584 l0bl12 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b12c585 l0bl12 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b12c586 l0bl12 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b12c587 l0bl12 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b12c588 l0bl12 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b12c589 l0bl12 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b12c590 l0bl12 vdd x590 x590b CELLD r1=10000e3 r0=900e3
xl0b12c591 l0bl12 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b12c592 l0bl12 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b12c593 l0bl12 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b12c594 l0bl12 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b12c595 l0bl12 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b12c596 l0bl12 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b12c597 l0bl12 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b12c598 l0bl12 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b12c599 l0bl12 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b12c600 l0bl12 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b12c601 l0bl12 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b12c602 l0bl12 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b12c603 l0bl12 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b12c604 l0bl12 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b12c605 l0bl12 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b12c606 l0bl12 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b12c607 l0bl12 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b12c608 l0bl12 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b12c609 l0bl12 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b12c610 l0bl12 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b12c611 l0bl12 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b12c612 l0bl12 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b12c613 l0bl12 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b12c614 l0bl12 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b12c615 l0bl12 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b12c616 l0bl12 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b12c617 l0bl12 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b12c618 l0bl12 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b12c619 l0bl12 vdd x619 x619b CELLD r1=900e3 r0=10000e3
xl0b12c620 l0bl12 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b12c621 l0bl12 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b12c622 l0bl12 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b12c623 l0bl12 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b12c624 l0bl12 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b12c625 l0bl12 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b12c626 l0bl12 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b12c627 l0bl12 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b12c628 l0bl12 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b12c629 l0bl12 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b12c630 l0bl12 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b12c631 l0bl12 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b12c632 l0bl12 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b12c633 l0bl12 vdd x633 x633b CELLD r1=10000e3 r0=900e3
xl0b12c634 l0bl12 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b12c635 l0bl12 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b12c636 l0bl12 vdd x636 x636b CELLD r1=10000e3 r0=900e3
xl0b12c637 l0bl12 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b12c638 l0bl12 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b12c639 l0bl12 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b12c640 l0bl12 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b12c641 l0bl12 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b12c642 l0bl12 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b12c643 l0bl12 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b12c644 l0bl12 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b12c645 l0bl12 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b12c646 l0bl12 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b12c647 l0bl12 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b12c648 l0bl12 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b12c649 l0bl12 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b12c650 l0bl12 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b12c651 l0bl12 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b12c652 l0bl12 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b12c653 l0bl12 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b12c654 l0bl12 vdd x654 x654b CELLD r1=900e3 r0=10000e3
xl0b12c655 l0bl12 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b12c656 l0bl12 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b12c657 l0bl12 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b12c658 l0bl12 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b12c659 l0bl12 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b12c660 l0bl12 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b12c661 l0bl12 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b12c662 l0bl12 vdd x662 x662b CELLD r1=10000e3 r0=900e3
xl0b12c663 l0bl12 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b12c664 l0bl12 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b12c665 l0bl12 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b12c666 l0bl12 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b12c667 l0bl12 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b12c668 l0bl12 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b12c669 l0bl12 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b12c670 l0bl12 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b12c671 l0bl12 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b12c672 l0bl12 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b12c673 l0bl12 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b12c674 l0bl12 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b12c675 l0bl12 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b12c676 l0bl12 vdd x676 x676b CELLD r1=900e3 r0=10000e3
xl0b12c677 l0bl12 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b12c678 l0bl12 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b12c679 l0bl12 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b12c680 l0bl12 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b12c681 l0bl12 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b12c682 l0bl12 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b12c683 l0bl12 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b12c684 l0bl12 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b12c685 l0bl12 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b12c686 l0bl12 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b12c687 l0bl12 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b12c688 l0bl12 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b12c689 l0bl12 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b12c690 l0bl12 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b12c691 l0bl12 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b12c692 l0bl12 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b12c693 l0bl12 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b12c694 l0bl12 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b12c695 l0bl12 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b12c696 l0bl12 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b12c697 l0bl12 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b12c698 l0bl12 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b12c699 l0bl12 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b12c700 l0bl12 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b12c701 l0bl12 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b12c702 l0bl12 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b12c703 l0bl12 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b12c704 l0bl12 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b12c705 l0bl12 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b12c706 l0bl12 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b12c707 l0bl12 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b12c708 l0bl12 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b12c709 l0bl12 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b12c710 l0bl12 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b12c711 l0bl12 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b12c712 l0bl12 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b12c713 l0bl12 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b12c714 l0bl12 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b12c715 l0bl12 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b12c716 l0bl12 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b12c717 l0bl12 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b12c718 l0bl12 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b12c719 l0bl12 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b12c720 l0bl12 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b12c721 l0bl12 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b12c722 l0bl12 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b12c723 l0bl12 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b12c724 l0bl12 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b12c725 l0bl12 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b12c726 l0bl12 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b12c727 l0bl12 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b12c728 l0bl12 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b12c729 l0bl12 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b12c730 l0bl12 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b12c731 l0bl12 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b12c732 l0bl12 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b12c733 l0bl12 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b12c734 l0bl12 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b12c735 l0bl12 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b12c736 l0bl12 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b12c737 l0bl12 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b12c738 l0bl12 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b12c739 l0bl12 vdd x739 x739b CELLD r1=900e3 r0=10000e3
xl0b12c740 l0bl12 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b12c741 l0bl12 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b12c742 l0bl12 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b12c743 l0bl12 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b12c744 l0bl12 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b12c745 l0bl12 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b12c746 l0bl12 vdd x746 x746b CELLD r1=900e3 r0=10000e3
xl0b12c747 l0bl12 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b12c748 l0bl12 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b12c749 l0bl12 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b12c750 l0bl12 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b12c751 l0bl12 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b12c752 l0bl12 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b12c753 l0bl12 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b12c754 l0bl12 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b12c755 l0bl12 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b12c756 l0bl12 vdd x756 x756b CELLD r1=900e3 r0=10000e3
xl0b12c757 l0bl12 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b12c758 l0bl12 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b12c759 l0bl12 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b12c760 l0bl12 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b12c761 l0bl12 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b12c762 l0bl12 vdd x762 x762b CELLD r1=900e3 r0=10000e3
xl0b12c763 l0bl12 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b12c764 l0bl12 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b12c765 l0bl12 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b12c766 l0bl12 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b12c767 l0bl12 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b12c768 l0bl12 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b12c769 l0bl12 vdd x769 x769b CELLD r1=900e3 r0=10000e3
xl0b12c770 l0bl12 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b12c771 l0bl12 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b12c772 l0bl12 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b12c773 l0bl12 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b12c774 l0bl12 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b12c775 l0bl12 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b12c776 l0bl12 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b12c777 l0bl12 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b12c778 l0bl12 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b12c779 l0bl12 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b12c780 l0bl12 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b12c781 l0bl12 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b12c782 l0bl12 vdd x782 x782b CELLD r1=10000e3 r0=900e3
xl0b12c783 l0bl12 vdd x783 x783b CELLD r1=900e3 r0=10000e3
xl0b13c0 l0bl13 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b13c1 l0bl13 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b13c2 l0bl13 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b13c3 l0bl13 vdd x3 x3b CELLD r1=10000e3 r0=900e3
xl0b13c4 l0bl13 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b13c5 l0bl13 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b13c6 l0bl13 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b13c7 l0bl13 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b13c8 l0bl13 vdd x8 x8b CELLD r1=900e3 r0=10000e3
xl0b13c9 l0bl13 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b13c10 l0bl13 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b13c11 l0bl13 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b13c12 l0bl13 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b13c13 l0bl13 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b13c14 l0bl13 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b13c15 l0bl13 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b13c16 l0bl13 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b13c17 l0bl13 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b13c18 l0bl13 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b13c19 l0bl13 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b13c20 l0bl13 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b13c21 l0bl13 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b13c22 l0bl13 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b13c23 l0bl13 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b13c24 l0bl13 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b13c25 l0bl13 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b13c26 l0bl13 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b13c27 l0bl13 vdd x27 x27b CELLD r1=900e3 r0=10000e3
xl0b13c28 l0bl13 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b13c29 l0bl13 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b13c30 l0bl13 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b13c31 l0bl13 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b13c32 l0bl13 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b13c33 l0bl13 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b13c34 l0bl13 vdd x34 x34b CELLD r1=10000e3 r0=900e3
xl0b13c35 l0bl13 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b13c36 l0bl13 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b13c37 l0bl13 vdd x37 x37b CELLD r1=900e3 r0=10000e3
xl0b13c38 l0bl13 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b13c39 l0bl13 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b13c40 l0bl13 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b13c41 l0bl13 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b13c42 l0bl13 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b13c43 l0bl13 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b13c44 l0bl13 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b13c45 l0bl13 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b13c46 l0bl13 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b13c47 l0bl13 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b13c48 l0bl13 vdd x48 x48b CELLD r1=900e3 r0=10000e3
xl0b13c49 l0bl13 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b13c50 l0bl13 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b13c51 l0bl13 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b13c52 l0bl13 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b13c53 l0bl13 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b13c54 l0bl13 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b13c55 l0bl13 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b13c56 l0bl13 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b13c57 l0bl13 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b13c58 l0bl13 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b13c59 l0bl13 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b13c60 l0bl13 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b13c61 l0bl13 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b13c62 l0bl13 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b13c63 l0bl13 vdd x63 x63b CELLD r1=900e3 r0=10000e3
xl0b13c64 l0bl13 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b13c65 l0bl13 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b13c66 l0bl13 vdd x66 x66b CELLD r1=900e3 r0=10000e3
xl0b13c67 l0bl13 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b13c68 l0bl13 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b13c69 l0bl13 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b13c70 l0bl13 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b13c71 l0bl13 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b13c72 l0bl13 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b13c73 l0bl13 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b13c74 l0bl13 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b13c75 l0bl13 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b13c76 l0bl13 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b13c77 l0bl13 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b13c78 l0bl13 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b13c79 l0bl13 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b13c80 l0bl13 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b13c81 l0bl13 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b13c82 l0bl13 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b13c83 l0bl13 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b13c84 l0bl13 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b13c85 l0bl13 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b13c86 l0bl13 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b13c87 l0bl13 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b13c88 l0bl13 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b13c89 l0bl13 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b13c90 l0bl13 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b13c91 l0bl13 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b13c92 l0bl13 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b13c93 l0bl13 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b13c94 l0bl13 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b13c95 l0bl13 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b13c96 l0bl13 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b13c97 l0bl13 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b13c98 l0bl13 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b13c99 l0bl13 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b13c100 l0bl13 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b13c101 l0bl13 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b13c102 l0bl13 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b13c103 l0bl13 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b13c104 l0bl13 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b13c105 l0bl13 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b13c106 l0bl13 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b13c107 l0bl13 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b13c108 l0bl13 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b13c109 l0bl13 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b13c110 l0bl13 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b13c111 l0bl13 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b13c112 l0bl13 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b13c113 l0bl13 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b13c114 l0bl13 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b13c115 l0bl13 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b13c116 l0bl13 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b13c117 l0bl13 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b13c118 l0bl13 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b13c119 l0bl13 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b13c120 l0bl13 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b13c121 l0bl13 vdd x121 x121b CELLD r1=900e3 r0=10000e3
xl0b13c122 l0bl13 vdd x122 x122b CELLD r1=900e3 r0=10000e3
xl0b13c123 l0bl13 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b13c124 l0bl13 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b13c125 l0bl13 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b13c126 l0bl13 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b13c127 l0bl13 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b13c128 l0bl13 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b13c129 l0bl13 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b13c130 l0bl13 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b13c131 l0bl13 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b13c132 l0bl13 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b13c133 l0bl13 vdd x133 x133b CELLD r1=10000e3 r0=900e3
xl0b13c134 l0bl13 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b13c135 l0bl13 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b13c136 l0bl13 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b13c137 l0bl13 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b13c138 l0bl13 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b13c139 l0bl13 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b13c140 l0bl13 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b13c141 l0bl13 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b13c142 l0bl13 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b13c143 l0bl13 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b13c144 l0bl13 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b13c145 l0bl13 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b13c146 l0bl13 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b13c147 l0bl13 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b13c148 l0bl13 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b13c149 l0bl13 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b13c150 l0bl13 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b13c151 l0bl13 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b13c152 l0bl13 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b13c153 l0bl13 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b13c154 l0bl13 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b13c155 l0bl13 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b13c156 l0bl13 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b13c157 l0bl13 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b13c158 l0bl13 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b13c159 l0bl13 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b13c160 l0bl13 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b13c161 l0bl13 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b13c162 l0bl13 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b13c163 l0bl13 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b13c164 l0bl13 vdd x164 x164b CELLD r1=10000e3 r0=900e3
xl0b13c165 l0bl13 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b13c166 l0bl13 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b13c167 l0bl13 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b13c168 l0bl13 vdd x168 x168b CELLD r1=900e3 r0=10000e3
xl0b13c169 l0bl13 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b13c170 l0bl13 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b13c171 l0bl13 vdd x171 x171b CELLD r1=10000e3 r0=900e3
xl0b13c172 l0bl13 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b13c173 l0bl13 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b13c174 l0bl13 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b13c175 l0bl13 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b13c176 l0bl13 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b13c177 l0bl13 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b13c178 l0bl13 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b13c179 l0bl13 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b13c180 l0bl13 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b13c181 l0bl13 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b13c182 l0bl13 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b13c183 l0bl13 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b13c184 l0bl13 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b13c185 l0bl13 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b13c186 l0bl13 vdd x186 x186b CELLD r1=10000e3 r0=900e3
xl0b13c187 l0bl13 vdd x187 x187b CELLD r1=10000e3 r0=900e3
xl0b13c188 l0bl13 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b13c189 l0bl13 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b13c190 l0bl13 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b13c191 l0bl13 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b13c192 l0bl13 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b13c193 l0bl13 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b13c194 l0bl13 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b13c195 l0bl13 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b13c196 l0bl13 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b13c197 l0bl13 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b13c198 l0bl13 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b13c199 l0bl13 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b13c200 l0bl13 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b13c201 l0bl13 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b13c202 l0bl13 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b13c203 l0bl13 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b13c204 l0bl13 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b13c205 l0bl13 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b13c206 l0bl13 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b13c207 l0bl13 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b13c208 l0bl13 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b13c209 l0bl13 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b13c210 l0bl13 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b13c211 l0bl13 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b13c212 l0bl13 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b13c213 l0bl13 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b13c214 l0bl13 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b13c215 l0bl13 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b13c216 l0bl13 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b13c217 l0bl13 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b13c218 l0bl13 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b13c219 l0bl13 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b13c220 l0bl13 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b13c221 l0bl13 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b13c222 l0bl13 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b13c223 l0bl13 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b13c224 l0bl13 vdd x224 x224b CELLD r1=900e3 r0=10000e3
xl0b13c225 l0bl13 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b13c226 l0bl13 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b13c227 l0bl13 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b13c228 l0bl13 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b13c229 l0bl13 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b13c230 l0bl13 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b13c231 l0bl13 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b13c232 l0bl13 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b13c233 l0bl13 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b13c234 l0bl13 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b13c235 l0bl13 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b13c236 l0bl13 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b13c237 l0bl13 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b13c238 l0bl13 vdd x238 x238b CELLD r1=10000e3 r0=900e3
xl0b13c239 l0bl13 vdd x239 x239b CELLD r1=10000e3 r0=900e3
xl0b13c240 l0bl13 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b13c241 l0bl13 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b13c242 l0bl13 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b13c243 l0bl13 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b13c244 l0bl13 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b13c245 l0bl13 vdd x245 x245b CELLD r1=900e3 r0=10000e3
xl0b13c246 l0bl13 vdd x246 x246b CELLD r1=900e3 r0=10000e3
xl0b13c247 l0bl13 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b13c248 l0bl13 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b13c249 l0bl13 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b13c250 l0bl13 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b13c251 l0bl13 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b13c252 l0bl13 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b13c253 l0bl13 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b13c254 l0bl13 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b13c255 l0bl13 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b13c256 l0bl13 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b13c257 l0bl13 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b13c258 l0bl13 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b13c259 l0bl13 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b13c260 l0bl13 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b13c261 l0bl13 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b13c262 l0bl13 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b13c263 l0bl13 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b13c264 l0bl13 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b13c265 l0bl13 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b13c266 l0bl13 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b13c267 l0bl13 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b13c268 l0bl13 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b13c269 l0bl13 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b13c270 l0bl13 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b13c271 l0bl13 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b13c272 l0bl13 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b13c273 l0bl13 vdd x273 x273b CELLD r1=900e3 r0=10000e3
xl0b13c274 l0bl13 vdd x274 x274b CELLD r1=900e3 r0=10000e3
xl0b13c275 l0bl13 vdd x275 x275b CELLD r1=900e3 r0=10000e3
xl0b13c276 l0bl13 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b13c277 l0bl13 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b13c278 l0bl13 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b13c279 l0bl13 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b13c280 l0bl13 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b13c281 l0bl13 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b13c282 l0bl13 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b13c283 l0bl13 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b13c284 l0bl13 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b13c285 l0bl13 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b13c286 l0bl13 vdd x286 x286b CELLD r1=900e3 r0=10000e3
xl0b13c287 l0bl13 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b13c288 l0bl13 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b13c289 l0bl13 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b13c290 l0bl13 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b13c291 l0bl13 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b13c292 l0bl13 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b13c293 l0bl13 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b13c294 l0bl13 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b13c295 l0bl13 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b13c296 l0bl13 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b13c297 l0bl13 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b13c298 l0bl13 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b13c299 l0bl13 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b13c300 l0bl13 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b13c301 l0bl13 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b13c302 l0bl13 vdd x302 x302b CELLD r1=900e3 r0=10000e3
xl0b13c303 l0bl13 vdd x303 x303b CELLD r1=900e3 r0=10000e3
xl0b13c304 l0bl13 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b13c305 l0bl13 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b13c306 l0bl13 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b13c307 l0bl13 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b13c308 l0bl13 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b13c309 l0bl13 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b13c310 l0bl13 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b13c311 l0bl13 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b13c312 l0bl13 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b13c313 l0bl13 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b13c314 l0bl13 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b13c315 l0bl13 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b13c316 l0bl13 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b13c317 l0bl13 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b13c318 l0bl13 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b13c319 l0bl13 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b13c320 l0bl13 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b13c321 l0bl13 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b13c322 l0bl13 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b13c323 l0bl13 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b13c324 l0bl13 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b13c325 l0bl13 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b13c326 l0bl13 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b13c327 l0bl13 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b13c328 l0bl13 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b13c329 l0bl13 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b13c330 l0bl13 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b13c331 l0bl13 vdd x331 x331b CELLD r1=900e3 r0=10000e3
xl0b13c332 l0bl13 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b13c333 l0bl13 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b13c334 l0bl13 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b13c335 l0bl13 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b13c336 l0bl13 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b13c337 l0bl13 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b13c338 l0bl13 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b13c339 l0bl13 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b13c340 l0bl13 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b13c341 l0bl13 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b13c342 l0bl13 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b13c343 l0bl13 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b13c344 l0bl13 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b13c345 l0bl13 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b13c346 l0bl13 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b13c347 l0bl13 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b13c348 l0bl13 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b13c349 l0bl13 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b13c350 l0bl13 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b13c351 l0bl13 vdd x351 x351b CELLD r1=10000e3 r0=900e3
xl0b13c352 l0bl13 vdd x352 x352b CELLD r1=10000e3 r0=900e3
xl0b13c353 l0bl13 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b13c354 l0bl13 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b13c355 l0bl13 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b13c356 l0bl13 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b13c357 l0bl13 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b13c358 l0bl13 vdd x358 x358b CELLD r1=900e3 r0=10000e3
xl0b13c359 l0bl13 vdd x359 x359b CELLD r1=900e3 r0=10000e3
xl0b13c360 l0bl13 vdd x360 x360b CELLD r1=900e3 r0=10000e3
xl0b13c361 l0bl13 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b13c362 l0bl13 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b13c363 l0bl13 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b13c364 l0bl13 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b13c365 l0bl13 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b13c366 l0bl13 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b13c367 l0bl13 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b13c368 l0bl13 vdd x368 x368b CELLD r1=900e3 r0=10000e3
xl0b13c369 l0bl13 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b13c370 l0bl13 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b13c371 l0bl13 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b13c372 l0bl13 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b13c373 l0bl13 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b13c374 l0bl13 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b13c375 l0bl13 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b13c376 l0bl13 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b13c377 l0bl13 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b13c378 l0bl13 vdd x378 x378b CELLD r1=10000e3 r0=900e3
xl0b13c379 l0bl13 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b13c380 l0bl13 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b13c381 l0bl13 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b13c382 l0bl13 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b13c383 l0bl13 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b13c384 l0bl13 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b13c385 l0bl13 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b13c386 l0bl13 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b13c387 l0bl13 vdd x387 x387b CELLD r1=900e3 r0=10000e3
xl0b13c388 l0bl13 vdd x388 x388b CELLD r1=900e3 r0=10000e3
xl0b13c389 l0bl13 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b13c390 l0bl13 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b13c391 l0bl13 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b13c392 l0bl13 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b13c393 l0bl13 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b13c394 l0bl13 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b13c395 l0bl13 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b13c396 l0bl13 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b13c397 l0bl13 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b13c398 l0bl13 vdd x398 x398b CELLD r1=900e3 r0=10000e3
xl0b13c399 l0bl13 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b13c400 l0bl13 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b13c401 l0bl13 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b13c402 l0bl13 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b13c403 l0bl13 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b13c404 l0bl13 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b13c405 l0bl13 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b13c406 l0bl13 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b13c407 l0bl13 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b13c408 l0bl13 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b13c409 l0bl13 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b13c410 l0bl13 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b13c411 l0bl13 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b13c412 l0bl13 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b13c413 l0bl13 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b13c414 l0bl13 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b13c415 l0bl13 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b13c416 l0bl13 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b13c417 l0bl13 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b13c418 l0bl13 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b13c419 l0bl13 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b13c420 l0bl13 vdd x420 x420b CELLD r1=10000e3 r0=900e3
xl0b13c421 l0bl13 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b13c422 l0bl13 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b13c423 l0bl13 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b13c424 l0bl13 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b13c425 l0bl13 vdd x425 x425b CELLD r1=900e3 r0=10000e3
xl0b13c426 l0bl13 vdd x426 x426b CELLD r1=900e3 r0=10000e3
xl0b13c427 l0bl13 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b13c428 l0bl13 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b13c429 l0bl13 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b13c430 l0bl13 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b13c431 l0bl13 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b13c432 l0bl13 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b13c433 l0bl13 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b13c434 l0bl13 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b13c435 l0bl13 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b13c436 l0bl13 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b13c437 l0bl13 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b13c438 l0bl13 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b13c439 l0bl13 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b13c440 l0bl13 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b13c441 l0bl13 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b13c442 l0bl13 vdd x442 x442b CELLD r1=900e3 r0=10000e3
xl0b13c443 l0bl13 vdd x443 x443b CELLD r1=900e3 r0=10000e3
xl0b13c444 l0bl13 vdd x444 x444b CELLD r1=900e3 r0=10000e3
xl0b13c445 l0bl13 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b13c446 l0bl13 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b13c447 l0bl13 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b13c448 l0bl13 vdd x448 x448b CELLD r1=10000e3 r0=900e3
xl0b13c449 l0bl13 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b13c450 l0bl13 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b13c451 l0bl13 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b13c452 l0bl13 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b13c453 l0bl13 vdd x453 x453b CELLD r1=900e3 r0=10000e3
xl0b13c454 l0bl13 vdd x454 x454b CELLD r1=900e3 r0=10000e3
xl0b13c455 l0bl13 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b13c456 l0bl13 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b13c457 l0bl13 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b13c458 l0bl13 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b13c459 l0bl13 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b13c460 l0bl13 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b13c461 l0bl13 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b13c462 l0bl13 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b13c463 l0bl13 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b13c464 l0bl13 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b13c465 l0bl13 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b13c466 l0bl13 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b13c467 l0bl13 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b13c468 l0bl13 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b13c469 l0bl13 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b13c470 l0bl13 vdd x470 x470b CELLD r1=900e3 r0=10000e3
xl0b13c471 l0bl13 vdd x471 x471b CELLD r1=900e3 r0=10000e3
xl0b13c472 l0bl13 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b13c473 l0bl13 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b13c474 l0bl13 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b13c475 l0bl13 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b13c476 l0bl13 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b13c477 l0bl13 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b13c478 l0bl13 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b13c479 l0bl13 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b13c480 l0bl13 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b13c481 l0bl13 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b13c482 l0bl13 vdd x482 x482b CELLD r1=900e3 r0=10000e3
xl0b13c483 l0bl13 vdd x483 x483b CELLD r1=900e3 r0=10000e3
xl0b13c484 l0bl13 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b13c485 l0bl13 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b13c486 l0bl13 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b13c487 l0bl13 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b13c488 l0bl13 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b13c489 l0bl13 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b13c490 l0bl13 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b13c491 l0bl13 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b13c492 l0bl13 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b13c493 l0bl13 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b13c494 l0bl13 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b13c495 l0bl13 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b13c496 l0bl13 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b13c497 l0bl13 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b13c498 l0bl13 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b13c499 l0bl13 vdd x499 x499b CELLD r1=900e3 r0=10000e3
xl0b13c500 l0bl13 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b13c501 l0bl13 vdd x501 x501b CELLD r1=900e3 r0=10000e3
xl0b13c502 l0bl13 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b13c503 l0bl13 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b13c504 l0bl13 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b13c505 l0bl13 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b13c506 l0bl13 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b13c507 l0bl13 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b13c508 l0bl13 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b13c509 l0bl13 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b13c510 l0bl13 vdd x510 x510b CELLD r1=900e3 r0=10000e3
xl0b13c511 l0bl13 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b13c512 l0bl13 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b13c513 l0bl13 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b13c514 l0bl13 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b13c515 l0bl13 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b13c516 l0bl13 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b13c517 l0bl13 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b13c518 l0bl13 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b13c519 l0bl13 vdd x519 x519b CELLD r1=900e3 r0=10000e3
xl0b13c520 l0bl13 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b13c521 l0bl13 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b13c522 l0bl13 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b13c523 l0bl13 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b13c524 l0bl13 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b13c525 l0bl13 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b13c526 l0bl13 vdd x526 x526b CELLD r1=900e3 r0=10000e3
xl0b13c527 l0bl13 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b13c528 l0bl13 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b13c529 l0bl13 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b13c530 l0bl13 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b13c531 l0bl13 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b13c532 l0bl13 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b13c533 l0bl13 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b13c534 l0bl13 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b13c535 l0bl13 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b13c536 l0bl13 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b13c537 l0bl13 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b13c538 l0bl13 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b13c539 l0bl13 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b13c540 l0bl13 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b13c541 l0bl13 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b13c542 l0bl13 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b13c543 l0bl13 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b13c544 l0bl13 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b13c545 l0bl13 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b13c546 l0bl13 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b13c547 l0bl13 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b13c548 l0bl13 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b13c549 l0bl13 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b13c550 l0bl13 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b13c551 l0bl13 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b13c552 l0bl13 vdd x552 x552b CELLD r1=900e3 r0=10000e3
xl0b13c553 l0bl13 vdd x553 x553b CELLD r1=900e3 r0=10000e3
xl0b13c554 l0bl13 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b13c555 l0bl13 vdd x555 x555b CELLD r1=900e3 r0=10000e3
xl0b13c556 l0bl13 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b13c557 l0bl13 vdd x557 x557b CELLD r1=900e3 r0=10000e3
xl0b13c558 l0bl13 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b13c559 l0bl13 vdd x559 x559b CELLD r1=900e3 r0=10000e3
xl0b13c560 l0bl13 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b13c561 l0bl13 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b13c562 l0bl13 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b13c563 l0bl13 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b13c564 l0bl13 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b13c565 l0bl13 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b13c566 l0bl13 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b13c567 l0bl13 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b13c568 l0bl13 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b13c569 l0bl13 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b13c570 l0bl13 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b13c571 l0bl13 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b13c572 l0bl13 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b13c573 l0bl13 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b13c574 l0bl13 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b13c575 l0bl13 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b13c576 l0bl13 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b13c577 l0bl13 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b13c578 l0bl13 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b13c579 l0bl13 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b13c580 l0bl13 vdd x580 x580b CELLD r1=900e3 r0=10000e3
xl0b13c581 l0bl13 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b13c582 l0bl13 vdd x582 x582b CELLD r1=900e3 r0=10000e3
xl0b13c583 l0bl13 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b13c584 l0bl13 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b13c585 l0bl13 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b13c586 l0bl13 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b13c587 l0bl13 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b13c588 l0bl13 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b13c589 l0bl13 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b13c590 l0bl13 vdd x590 x590b CELLD r1=10000e3 r0=900e3
xl0b13c591 l0bl13 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b13c592 l0bl13 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b13c593 l0bl13 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b13c594 l0bl13 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b13c595 l0bl13 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b13c596 l0bl13 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b13c597 l0bl13 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b13c598 l0bl13 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b13c599 l0bl13 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b13c600 l0bl13 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b13c601 l0bl13 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b13c602 l0bl13 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b13c603 l0bl13 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b13c604 l0bl13 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b13c605 l0bl13 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b13c606 l0bl13 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b13c607 l0bl13 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b13c608 l0bl13 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b13c609 l0bl13 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b13c610 l0bl13 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b13c611 l0bl13 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b13c612 l0bl13 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b13c613 l0bl13 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b13c614 l0bl13 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b13c615 l0bl13 vdd x615 x615b CELLD r1=900e3 r0=10000e3
xl0b13c616 l0bl13 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b13c617 l0bl13 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b13c618 l0bl13 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b13c619 l0bl13 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b13c620 l0bl13 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b13c621 l0bl13 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b13c622 l0bl13 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b13c623 l0bl13 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b13c624 l0bl13 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b13c625 l0bl13 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b13c626 l0bl13 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b13c627 l0bl13 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b13c628 l0bl13 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b13c629 l0bl13 vdd x629 x629b CELLD r1=900e3 r0=10000e3
xl0b13c630 l0bl13 vdd x630 x630b CELLD r1=900e3 r0=10000e3
xl0b13c631 l0bl13 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b13c632 l0bl13 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b13c633 l0bl13 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b13c634 l0bl13 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b13c635 l0bl13 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b13c636 l0bl13 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b13c637 l0bl13 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b13c638 l0bl13 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b13c639 l0bl13 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b13c640 l0bl13 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b13c641 l0bl13 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b13c642 l0bl13 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b13c643 l0bl13 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b13c644 l0bl13 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b13c645 l0bl13 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b13c646 l0bl13 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b13c647 l0bl13 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b13c648 l0bl13 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b13c649 l0bl13 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b13c650 l0bl13 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b13c651 l0bl13 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b13c652 l0bl13 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b13c653 l0bl13 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b13c654 l0bl13 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b13c655 l0bl13 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b13c656 l0bl13 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b13c657 l0bl13 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b13c658 l0bl13 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b13c659 l0bl13 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b13c660 l0bl13 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b13c661 l0bl13 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b13c662 l0bl13 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b13c663 l0bl13 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b13c664 l0bl13 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b13c665 l0bl13 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b13c666 l0bl13 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b13c667 l0bl13 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b13c668 l0bl13 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b13c669 l0bl13 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b13c670 l0bl13 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b13c671 l0bl13 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b13c672 l0bl13 vdd x672 x672b CELLD r1=900e3 r0=10000e3
xl0b13c673 l0bl13 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b13c674 l0bl13 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b13c675 l0bl13 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b13c676 l0bl13 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b13c677 l0bl13 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b13c678 l0bl13 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b13c679 l0bl13 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b13c680 l0bl13 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b13c681 l0bl13 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b13c682 l0bl13 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b13c683 l0bl13 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b13c684 l0bl13 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b13c685 l0bl13 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b13c686 l0bl13 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b13c687 l0bl13 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b13c688 l0bl13 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b13c689 l0bl13 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b13c690 l0bl13 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b13c691 l0bl13 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b13c692 l0bl13 vdd x692 x692b CELLD r1=10000e3 r0=900e3
xl0b13c693 l0bl13 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b13c694 l0bl13 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b13c695 l0bl13 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b13c696 l0bl13 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b13c697 l0bl13 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b13c698 l0bl13 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b13c699 l0bl13 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b13c700 l0bl13 vdd x700 x700b CELLD r1=900e3 r0=10000e3
xl0b13c701 l0bl13 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b13c702 l0bl13 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b13c703 l0bl13 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b13c704 l0bl13 vdd x704 x704b CELLD r1=10000e3 r0=900e3
xl0b13c705 l0bl13 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b13c706 l0bl13 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b13c707 l0bl13 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b13c708 l0bl13 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b13c709 l0bl13 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b13c710 l0bl13 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b13c711 l0bl13 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b13c712 l0bl13 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b13c713 l0bl13 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b13c714 l0bl13 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b13c715 l0bl13 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b13c716 l0bl13 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b13c717 l0bl13 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b13c718 l0bl13 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b13c719 l0bl13 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b13c720 l0bl13 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b13c721 l0bl13 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b13c722 l0bl13 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b13c723 l0bl13 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b13c724 l0bl13 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b13c725 l0bl13 vdd x725 x725b CELLD r1=10000e3 r0=900e3
xl0b13c726 l0bl13 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b13c727 l0bl13 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b13c728 l0bl13 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b13c729 l0bl13 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b13c730 l0bl13 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b13c731 l0bl13 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b13c732 l0bl13 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b13c733 l0bl13 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b13c734 l0bl13 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b13c735 l0bl13 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b13c736 l0bl13 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b13c737 l0bl13 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b13c738 l0bl13 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b13c739 l0bl13 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b13c740 l0bl13 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b13c741 l0bl13 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b13c742 l0bl13 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b13c743 l0bl13 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b13c744 l0bl13 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b13c745 l0bl13 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b13c746 l0bl13 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b13c747 l0bl13 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b13c748 l0bl13 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b13c749 l0bl13 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b13c750 l0bl13 vdd x750 x750b CELLD r1=10000e3 r0=900e3
xl0b13c751 l0bl13 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b13c752 l0bl13 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b13c753 l0bl13 vdd x753 x753b CELLD r1=900e3 r0=10000e3
xl0b13c754 l0bl13 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b13c755 l0bl13 vdd x755 x755b CELLD r1=10000e3 r0=900e3
xl0b13c756 l0bl13 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b13c757 l0bl13 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b13c758 l0bl13 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b13c759 l0bl13 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b13c760 l0bl13 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b13c761 l0bl13 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b13c762 l0bl13 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b13c763 l0bl13 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b13c764 l0bl13 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b13c765 l0bl13 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b13c766 l0bl13 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b13c767 l0bl13 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b13c768 l0bl13 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b13c769 l0bl13 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b13c770 l0bl13 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b13c771 l0bl13 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b13c772 l0bl13 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b13c773 l0bl13 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b13c774 l0bl13 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b13c775 l0bl13 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b13c776 l0bl13 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b13c777 l0bl13 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b13c778 l0bl13 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b13c779 l0bl13 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b13c780 l0bl13 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b13c781 l0bl13 vdd x781 x781b CELLD r1=10000e3 r0=900e3
xl0b13c782 l0bl13 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b13c783 l0bl13 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b14c0 l0bl14 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b14c1 l0bl14 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b14c2 l0bl14 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b14c3 l0bl14 vdd x3 x3b CELLD r1=10000e3 r0=900e3
xl0b14c4 l0bl14 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b14c5 l0bl14 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b14c6 l0bl14 vdd x6 x6b CELLD r1=10000e3 r0=900e3
xl0b14c7 l0bl14 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b14c8 l0bl14 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b14c9 l0bl14 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b14c10 l0bl14 vdd x10 x10b CELLD r1=10000e3 r0=900e3
xl0b14c11 l0bl14 vdd x11 x11b CELLD r1=10000e3 r0=900e3
xl0b14c12 l0bl14 vdd x12 x12b CELLD r1=10000e3 r0=900e3
xl0b14c13 l0bl14 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b14c14 l0bl14 vdd x14 x14b CELLD r1=10000e3 r0=900e3
xl0b14c15 l0bl14 vdd x15 x15b CELLD r1=10000e3 r0=900e3
xl0b14c16 l0bl14 vdd x16 x16b CELLD r1=10000e3 r0=900e3
xl0b14c17 l0bl14 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b14c18 l0bl14 vdd x18 x18b CELLD r1=10000e3 r0=900e3
xl0b14c19 l0bl14 vdd x19 x19b CELLD r1=10000e3 r0=900e3
xl0b14c20 l0bl14 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b14c21 l0bl14 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b14c22 l0bl14 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b14c23 l0bl14 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b14c24 l0bl14 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b14c25 l0bl14 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b14c26 l0bl14 vdd x26 x26b CELLD r1=10000e3 r0=900e3
xl0b14c27 l0bl14 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b14c28 l0bl14 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b14c29 l0bl14 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b14c30 l0bl14 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b14c31 l0bl14 vdd x31 x31b CELLD r1=10000e3 r0=900e3
xl0b14c32 l0bl14 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b14c33 l0bl14 vdd x33 x33b CELLD r1=10000e3 r0=900e3
xl0b14c34 l0bl14 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b14c35 l0bl14 vdd x35 x35b CELLD r1=10000e3 r0=900e3
xl0b14c36 l0bl14 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b14c37 l0bl14 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b14c38 l0bl14 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b14c39 l0bl14 vdd x39 x39b CELLD r1=10000e3 r0=900e3
xl0b14c40 l0bl14 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b14c41 l0bl14 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b14c42 l0bl14 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b14c43 l0bl14 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b14c44 l0bl14 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b14c45 l0bl14 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b14c46 l0bl14 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b14c47 l0bl14 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b14c48 l0bl14 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b14c49 l0bl14 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b14c50 l0bl14 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b14c51 l0bl14 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b14c52 l0bl14 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b14c53 l0bl14 vdd x53 x53b CELLD r1=900e3 r0=10000e3
xl0b14c54 l0bl14 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b14c55 l0bl14 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b14c56 l0bl14 vdd x56 x56b CELLD r1=10000e3 r0=900e3
xl0b14c57 l0bl14 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b14c58 l0bl14 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b14c59 l0bl14 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b14c60 l0bl14 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b14c61 l0bl14 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b14c62 l0bl14 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b14c63 l0bl14 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b14c64 l0bl14 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b14c65 l0bl14 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b14c66 l0bl14 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b14c67 l0bl14 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b14c68 l0bl14 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b14c69 l0bl14 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b14c70 l0bl14 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b14c71 l0bl14 vdd x71 x71b CELLD r1=900e3 r0=10000e3
xl0b14c72 l0bl14 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b14c73 l0bl14 vdd x73 x73b CELLD r1=900e3 r0=10000e3
xl0b14c74 l0bl14 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b14c75 l0bl14 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b14c76 l0bl14 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b14c77 l0bl14 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b14c78 l0bl14 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b14c79 l0bl14 vdd x79 x79b CELLD r1=10000e3 r0=900e3
xl0b14c80 l0bl14 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b14c81 l0bl14 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b14c82 l0bl14 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b14c83 l0bl14 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b14c84 l0bl14 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b14c85 l0bl14 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b14c86 l0bl14 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b14c87 l0bl14 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b14c88 l0bl14 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b14c89 l0bl14 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b14c90 l0bl14 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b14c91 l0bl14 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b14c92 l0bl14 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b14c93 l0bl14 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b14c94 l0bl14 vdd x94 x94b CELLD r1=900e3 r0=10000e3
xl0b14c95 l0bl14 vdd x95 x95b CELLD r1=900e3 r0=10000e3
xl0b14c96 l0bl14 vdd x96 x96b CELLD r1=900e3 r0=10000e3
xl0b14c97 l0bl14 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b14c98 l0bl14 vdd x98 x98b CELLD r1=900e3 r0=10000e3
xl0b14c99 l0bl14 vdd x99 x99b CELLD r1=900e3 r0=10000e3
xl0b14c100 l0bl14 vdd x100 x100b CELLD r1=900e3 r0=10000e3
xl0b14c101 l0bl14 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b14c102 l0bl14 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b14c103 l0bl14 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b14c104 l0bl14 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b14c105 l0bl14 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b14c106 l0bl14 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b14c107 l0bl14 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b14c108 l0bl14 vdd x108 x108b CELLD r1=10000e3 r0=900e3
xl0b14c109 l0bl14 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b14c110 l0bl14 vdd x110 x110b CELLD r1=10000e3 r0=900e3
xl0b14c111 l0bl14 vdd x111 x111b CELLD r1=10000e3 r0=900e3
xl0b14c112 l0bl14 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b14c113 l0bl14 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b14c114 l0bl14 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b14c115 l0bl14 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b14c116 l0bl14 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b14c117 l0bl14 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b14c118 l0bl14 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b14c119 l0bl14 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b14c120 l0bl14 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b14c121 l0bl14 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b14c122 l0bl14 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b14c123 l0bl14 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b14c124 l0bl14 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b14c125 l0bl14 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b14c126 l0bl14 vdd x126 x126b CELLD r1=900e3 r0=10000e3
xl0b14c127 l0bl14 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b14c128 l0bl14 vdd x128 x128b CELLD r1=900e3 r0=10000e3
xl0b14c129 l0bl14 vdd x129 x129b CELLD r1=900e3 r0=10000e3
xl0b14c130 l0bl14 vdd x130 x130b CELLD r1=900e3 r0=10000e3
xl0b14c131 l0bl14 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b14c132 l0bl14 vdd x132 x132b CELLD r1=10000e3 r0=900e3
xl0b14c133 l0bl14 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b14c134 l0bl14 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b14c135 l0bl14 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b14c136 l0bl14 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b14c137 l0bl14 vdd x137 x137b CELLD r1=10000e3 r0=900e3
xl0b14c138 l0bl14 vdd x138 x138b CELLD r1=10000e3 r0=900e3
xl0b14c139 l0bl14 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b14c140 l0bl14 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b14c141 l0bl14 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b14c142 l0bl14 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b14c143 l0bl14 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b14c144 l0bl14 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b14c145 l0bl14 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b14c146 l0bl14 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b14c147 l0bl14 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b14c148 l0bl14 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b14c149 l0bl14 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b14c150 l0bl14 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b14c151 l0bl14 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b14c152 l0bl14 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b14c153 l0bl14 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b14c154 l0bl14 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b14c155 l0bl14 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b14c156 l0bl14 vdd x156 x156b CELLD r1=900e3 r0=10000e3
xl0b14c157 l0bl14 vdd x157 x157b CELLD r1=900e3 r0=10000e3
xl0b14c158 l0bl14 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b14c159 l0bl14 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b14c160 l0bl14 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b14c161 l0bl14 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b14c162 l0bl14 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b14c163 l0bl14 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b14c164 l0bl14 vdd x164 x164b CELLD r1=10000e3 r0=900e3
xl0b14c165 l0bl14 vdd x165 x165b CELLD r1=10000e3 r0=900e3
xl0b14c166 l0bl14 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b14c167 l0bl14 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b14c168 l0bl14 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b14c169 l0bl14 vdd x169 x169b CELLD r1=10000e3 r0=900e3
xl0b14c170 l0bl14 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b14c171 l0bl14 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b14c172 l0bl14 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b14c173 l0bl14 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b14c174 l0bl14 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b14c175 l0bl14 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b14c176 l0bl14 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b14c177 l0bl14 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b14c178 l0bl14 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b14c179 l0bl14 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b14c180 l0bl14 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b14c181 l0bl14 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b14c182 l0bl14 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b14c183 l0bl14 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b14c184 l0bl14 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b14c185 l0bl14 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b14c186 l0bl14 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b14c187 l0bl14 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b14c188 l0bl14 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b14c189 l0bl14 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b14c190 l0bl14 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b14c191 l0bl14 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b14c192 l0bl14 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b14c193 l0bl14 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b14c194 l0bl14 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b14c195 l0bl14 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b14c196 l0bl14 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b14c197 l0bl14 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b14c198 l0bl14 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b14c199 l0bl14 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b14c200 l0bl14 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b14c201 l0bl14 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b14c202 l0bl14 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b14c203 l0bl14 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b14c204 l0bl14 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b14c205 l0bl14 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b14c206 l0bl14 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b14c207 l0bl14 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b14c208 l0bl14 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b14c209 l0bl14 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b14c210 l0bl14 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b14c211 l0bl14 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b14c212 l0bl14 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b14c213 l0bl14 vdd x213 x213b CELLD r1=10000e3 r0=900e3
xl0b14c214 l0bl14 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b14c215 l0bl14 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b14c216 l0bl14 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b14c217 l0bl14 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b14c218 l0bl14 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b14c219 l0bl14 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b14c220 l0bl14 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b14c221 l0bl14 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b14c222 l0bl14 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b14c223 l0bl14 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b14c224 l0bl14 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b14c225 l0bl14 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b14c226 l0bl14 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b14c227 l0bl14 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b14c228 l0bl14 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b14c229 l0bl14 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b14c230 l0bl14 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b14c231 l0bl14 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b14c232 l0bl14 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b14c233 l0bl14 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b14c234 l0bl14 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b14c235 l0bl14 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b14c236 l0bl14 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b14c237 l0bl14 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b14c238 l0bl14 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b14c239 l0bl14 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b14c240 l0bl14 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b14c241 l0bl14 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b14c242 l0bl14 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b14c243 l0bl14 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b14c244 l0bl14 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b14c245 l0bl14 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b14c246 l0bl14 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b14c247 l0bl14 vdd x247 x247b CELLD r1=900e3 r0=10000e3
xl0b14c248 l0bl14 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b14c249 l0bl14 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b14c250 l0bl14 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b14c251 l0bl14 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b14c252 l0bl14 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b14c253 l0bl14 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b14c254 l0bl14 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b14c255 l0bl14 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b14c256 l0bl14 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b14c257 l0bl14 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b14c258 l0bl14 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b14c259 l0bl14 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b14c260 l0bl14 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b14c261 l0bl14 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b14c262 l0bl14 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b14c263 l0bl14 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b14c264 l0bl14 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b14c265 l0bl14 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b14c266 l0bl14 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b14c267 l0bl14 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b14c268 l0bl14 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b14c269 l0bl14 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b14c270 l0bl14 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b14c271 l0bl14 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b14c272 l0bl14 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b14c273 l0bl14 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b14c274 l0bl14 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b14c275 l0bl14 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b14c276 l0bl14 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b14c277 l0bl14 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b14c278 l0bl14 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b14c279 l0bl14 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b14c280 l0bl14 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b14c281 l0bl14 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b14c282 l0bl14 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b14c283 l0bl14 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b14c284 l0bl14 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b14c285 l0bl14 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b14c286 l0bl14 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b14c287 l0bl14 vdd x287 x287b CELLD r1=900e3 r0=10000e3
xl0b14c288 l0bl14 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b14c289 l0bl14 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b14c290 l0bl14 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b14c291 l0bl14 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b14c292 l0bl14 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b14c293 l0bl14 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b14c294 l0bl14 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b14c295 l0bl14 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b14c296 l0bl14 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b14c297 l0bl14 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b14c298 l0bl14 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b14c299 l0bl14 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b14c300 l0bl14 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b14c301 l0bl14 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b14c302 l0bl14 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b14c303 l0bl14 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b14c304 l0bl14 vdd x304 x304b CELLD r1=900e3 r0=10000e3
xl0b14c305 l0bl14 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b14c306 l0bl14 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b14c307 l0bl14 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b14c308 l0bl14 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b14c309 l0bl14 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b14c310 l0bl14 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b14c311 l0bl14 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b14c312 l0bl14 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b14c313 l0bl14 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b14c314 l0bl14 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b14c315 l0bl14 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b14c316 l0bl14 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b14c317 l0bl14 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b14c318 l0bl14 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b14c319 l0bl14 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b14c320 l0bl14 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b14c321 l0bl14 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b14c322 l0bl14 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b14c323 l0bl14 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b14c324 l0bl14 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b14c325 l0bl14 vdd x325 x325b CELLD r1=10000e3 r0=900e3
xl0b14c326 l0bl14 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b14c327 l0bl14 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b14c328 l0bl14 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b14c329 l0bl14 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b14c330 l0bl14 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b14c331 l0bl14 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b14c332 l0bl14 vdd x332 x332b CELLD r1=900e3 r0=10000e3
xl0b14c333 l0bl14 vdd x333 x333b CELLD r1=900e3 r0=10000e3
xl0b14c334 l0bl14 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b14c335 l0bl14 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b14c336 l0bl14 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b14c337 l0bl14 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b14c338 l0bl14 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b14c339 l0bl14 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b14c340 l0bl14 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b14c341 l0bl14 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b14c342 l0bl14 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b14c343 l0bl14 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b14c344 l0bl14 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b14c345 l0bl14 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b14c346 l0bl14 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b14c347 l0bl14 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b14c348 l0bl14 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b14c349 l0bl14 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b14c350 l0bl14 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b14c351 l0bl14 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b14c352 l0bl14 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b14c353 l0bl14 vdd x353 x353b CELLD r1=10000e3 r0=900e3
xl0b14c354 l0bl14 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b14c355 l0bl14 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b14c356 l0bl14 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b14c357 l0bl14 vdd x357 x357b CELLD r1=900e3 r0=10000e3
xl0b14c358 l0bl14 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b14c359 l0bl14 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b14c360 l0bl14 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b14c361 l0bl14 vdd x361 x361b CELLD r1=900e3 r0=10000e3
xl0b14c362 l0bl14 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b14c363 l0bl14 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b14c364 l0bl14 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b14c365 l0bl14 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b14c366 l0bl14 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b14c367 l0bl14 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b14c368 l0bl14 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b14c369 l0bl14 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b14c370 l0bl14 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b14c371 l0bl14 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b14c372 l0bl14 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b14c373 l0bl14 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b14c374 l0bl14 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b14c375 l0bl14 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b14c376 l0bl14 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b14c377 l0bl14 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b14c378 l0bl14 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b14c379 l0bl14 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b14c380 l0bl14 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b14c381 l0bl14 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b14c382 l0bl14 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b14c383 l0bl14 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b14c384 l0bl14 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b14c385 l0bl14 vdd x385 x385b CELLD r1=900e3 r0=10000e3
xl0b14c386 l0bl14 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b14c387 l0bl14 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b14c388 l0bl14 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b14c389 l0bl14 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b14c390 l0bl14 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b14c391 l0bl14 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b14c392 l0bl14 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b14c393 l0bl14 vdd x393 x393b CELLD r1=10000e3 r0=900e3
xl0b14c394 l0bl14 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b14c395 l0bl14 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b14c396 l0bl14 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b14c397 l0bl14 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b14c398 l0bl14 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b14c399 l0bl14 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b14c400 l0bl14 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b14c401 l0bl14 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b14c402 l0bl14 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b14c403 l0bl14 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b14c404 l0bl14 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b14c405 l0bl14 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b14c406 l0bl14 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b14c407 l0bl14 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b14c408 l0bl14 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b14c409 l0bl14 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b14c410 l0bl14 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b14c411 l0bl14 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b14c412 l0bl14 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b14c413 l0bl14 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b14c414 l0bl14 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b14c415 l0bl14 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b14c416 l0bl14 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b14c417 l0bl14 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b14c418 l0bl14 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b14c419 l0bl14 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b14c420 l0bl14 vdd x420 x420b CELLD r1=10000e3 r0=900e3
xl0b14c421 l0bl14 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b14c422 l0bl14 vdd x422 x422b CELLD r1=10000e3 r0=900e3
xl0b14c423 l0bl14 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b14c424 l0bl14 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b14c425 l0bl14 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b14c426 l0bl14 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b14c427 l0bl14 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b14c428 l0bl14 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b14c429 l0bl14 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b14c430 l0bl14 vdd x430 x430b CELLD r1=10000e3 r0=900e3
xl0b14c431 l0bl14 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b14c432 l0bl14 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b14c433 l0bl14 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b14c434 l0bl14 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b14c435 l0bl14 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b14c436 l0bl14 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b14c437 l0bl14 vdd x437 x437b CELLD r1=10000e3 r0=900e3
xl0b14c438 l0bl14 vdd x438 x438b CELLD r1=10000e3 r0=900e3
xl0b14c439 l0bl14 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b14c440 l0bl14 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b14c441 l0bl14 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b14c442 l0bl14 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b14c443 l0bl14 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b14c444 l0bl14 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b14c445 l0bl14 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b14c446 l0bl14 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b14c447 l0bl14 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b14c448 l0bl14 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b14c449 l0bl14 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b14c450 l0bl14 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b14c451 l0bl14 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b14c452 l0bl14 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b14c453 l0bl14 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b14c454 l0bl14 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b14c455 l0bl14 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b14c456 l0bl14 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b14c457 l0bl14 vdd x457 x457b CELLD r1=10000e3 r0=900e3
xl0b14c458 l0bl14 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b14c459 l0bl14 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b14c460 l0bl14 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b14c461 l0bl14 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b14c462 l0bl14 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b14c463 l0bl14 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b14c464 l0bl14 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b14c465 l0bl14 vdd x465 x465b CELLD r1=10000e3 r0=900e3
xl0b14c466 l0bl14 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b14c467 l0bl14 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b14c468 l0bl14 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b14c469 l0bl14 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b14c470 l0bl14 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b14c471 l0bl14 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b14c472 l0bl14 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b14c473 l0bl14 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b14c474 l0bl14 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b14c475 l0bl14 vdd x475 x475b CELLD r1=10000e3 r0=900e3
xl0b14c476 l0bl14 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b14c477 l0bl14 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b14c478 l0bl14 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b14c479 l0bl14 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b14c480 l0bl14 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b14c481 l0bl14 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b14c482 l0bl14 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b14c483 l0bl14 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b14c484 l0bl14 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b14c485 l0bl14 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b14c486 l0bl14 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b14c487 l0bl14 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b14c488 l0bl14 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b14c489 l0bl14 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b14c490 l0bl14 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b14c491 l0bl14 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b14c492 l0bl14 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b14c493 l0bl14 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b14c494 l0bl14 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b14c495 l0bl14 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b14c496 l0bl14 vdd x496 x496b CELLD r1=900e3 r0=10000e3
xl0b14c497 l0bl14 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b14c498 l0bl14 vdd x498 x498b CELLD r1=900e3 r0=10000e3
xl0b14c499 l0bl14 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b14c500 l0bl14 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b14c501 l0bl14 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b14c502 l0bl14 vdd x502 x502b CELLD r1=900e3 r0=10000e3
xl0b14c503 l0bl14 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b14c504 l0bl14 vdd x504 x504b CELLD r1=10000e3 r0=900e3
xl0b14c505 l0bl14 vdd x505 x505b CELLD r1=10000e3 r0=900e3
xl0b14c506 l0bl14 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b14c507 l0bl14 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b14c508 l0bl14 vdd x508 x508b CELLD r1=900e3 r0=10000e3
xl0b14c509 l0bl14 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b14c510 l0bl14 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b14c511 l0bl14 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b14c512 l0bl14 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b14c513 l0bl14 vdd x513 x513b CELLD r1=10000e3 r0=900e3
xl0b14c514 l0bl14 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b14c515 l0bl14 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b14c516 l0bl14 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b14c517 l0bl14 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b14c518 l0bl14 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b14c519 l0bl14 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b14c520 l0bl14 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b14c521 l0bl14 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b14c522 l0bl14 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b14c523 l0bl14 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b14c524 l0bl14 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b14c525 l0bl14 vdd x525 x525b CELLD r1=900e3 r0=10000e3
xl0b14c526 l0bl14 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b14c527 l0bl14 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b14c528 l0bl14 vdd x528 x528b CELLD r1=900e3 r0=10000e3
xl0b14c529 l0bl14 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b14c530 l0bl14 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b14c531 l0bl14 vdd x531 x531b CELLD r1=10000e3 r0=900e3
xl0b14c532 l0bl14 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b14c533 l0bl14 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b14c534 l0bl14 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b14c535 l0bl14 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b14c536 l0bl14 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b14c537 l0bl14 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b14c538 l0bl14 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b14c539 l0bl14 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b14c540 l0bl14 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b14c541 l0bl14 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b14c542 l0bl14 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b14c543 l0bl14 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b14c544 l0bl14 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b14c545 l0bl14 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b14c546 l0bl14 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b14c547 l0bl14 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b14c548 l0bl14 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b14c549 l0bl14 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b14c550 l0bl14 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b14c551 l0bl14 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b14c552 l0bl14 vdd x552 x552b CELLD r1=900e3 r0=10000e3
xl0b14c553 l0bl14 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b14c554 l0bl14 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b14c555 l0bl14 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b14c556 l0bl14 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b14c557 l0bl14 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b14c558 l0bl14 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b14c559 l0bl14 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b14c560 l0bl14 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b14c561 l0bl14 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b14c562 l0bl14 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b14c563 l0bl14 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b14c564 l0bl14 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b14c565 l0bl14 vdd x565 x565b CELLD r1=900e3 r0=10000e3
xl0b14c566 l0bl14 vdd x566 x566b CELLD r1=900e3 r0=10000e3
xl0b14c567 l0bl14 vdd x567 x567b CELLD r1=900e3 r0=10000e3
xl0b14c568 l0bl14 vdd x568 x568b CELLD r1=900e3 r0=10000e3
xl0b14c569 l0bl14 vdd x569 x569b CELLD r1=900e3 r0=10000e3
xl0b14c570 l0bl14 vdd x570 x570b CELLD r1=900e3 r0=10000e3
xl0b14c571 l0bl14 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b14c572 l0bl14 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b14c573 l0bl14 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b14c574 l0bl14 vdd x574 x574b CELLD r1=900e3 r0=10000e3
xl0b14c575 l0bl14 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b14c576 l0bl14 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b14c577 l0bl14 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b14c578 l0bl14 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b14c579 l0bl14 vdd x579 x579b CELLD r1=900e3 r0=10000e3
xl0b14c580 l0bl14 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b14c581 l0bl14 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b14c582 l0bl14 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b14c583 l0bl14 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b14c584 l0bl14 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b14c585 l0bl14 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b14c586 l0bl14 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b14c587 l0bl14 vdd x587 x587b CELLD r1=10000e3 r0=900e3
xl0b14c588 l0bl14 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b14c589 l0bl14 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b14c590 l0bl14 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b14c591 l0bl14 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b14c592 l0bl14 vdd x592 x592b CELLD r1=900e3 r0=10000e3
xl0b14c593 l0bl14 vdd x593 x593b CELLD r1=900e3 r0=10000e3
xl0b14c594 l0bl14 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b14c595 l0bl14 vdd x595 x595b CELLD r1=900e3 r0=10000e3
xl0b14c596 l0bl14 vdd x596 x596b CELLD r1=900e3 r0=10000e3
xl0b14c597 l0bl14 vdd x597 x597b CELLD r1=900e3 r0=10000e3
xl0b14c598 l0bl14 vdd x598 x598b CELLD r1=900e3 r0=10000e3
xl0b14c599 l0bl14 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b14c600 l0bl14 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b14c601 l0bl14 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b14c602 l0bl14 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b14c603 l0bl14 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b14c604 l0bl14 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b14c605 l0bl14 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b14c606 l0bl14 vdd x606 x606b CELLD r1=900e3 r0=10000e3
xl0b14c607 l0bl14 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b14c608 l0bl14 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b14c609 l0bl14 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b14c610 l0bl14 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b14c611 l0bl14 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b14c612 l0bl14 vdd x612 x612b CELLD r1=900e3 r0=10000e3
xl0b14c613 l0bl14 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b14c614 l0bl14 vdd x614 x614b CELLD r1=10000e3 r0=900e3
xl0b14c615 l0bl14 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b14c616 l0bl14 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b14c617 l0bl14 vdd x617 x617b CELLD r1=10000e3 r0=900e3
xl0b14c618 l0bl14 vdd x618 x618b CELLD r1=10000e3 r0=900e3
xl0b14c619 l0bl14 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b14c620 l0bl14 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b14c621 l0bl14 vdd x621 x621b CELLD r1=900e3 r0=10000e3
xl0b14c622 l0bl14 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b14c623 l0bl14 vdd x623 x623b CELLD r1=900e3 r0=10000e3
xl0b14c624 l0bl14 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b14c625 l0bl14 vdd x625 x625b CELLD r1=900e3 r0=10000e3
xl0b14c626 l0bl14 vdd x626 x626b CELLD r1=900e3 r0=10000e3
xl0b14c627 l0bl14 vdd x627 x627b CELLD r1=900e3 r0=10000e3
xl0b14c628 l0bl14 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b14c629 l0bl14 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b14c630 l0bl14 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b14c631 l0bl14 vdd x631 x631b CELLD r1=900e3 r0=10000e3
xl0b14c632 l0bl14 vdd x632 x632b CELLD r1=900e3 r0=10000e3
xl0b14c633 l0bl14 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b14c634 l0bl14 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b14c635 l0bl14 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b14c636 l0bl14 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b14c637 l0bl14 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b14c638 l0bl14 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b14c639 l0bl14 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b14c640 l0bl14 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b14c641 l0bl14 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b14c642 l0bl14 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b14c643 l0bl14 vdd x643 x643b CELLD r1=10000e3 r0=900e3
xl0b14c644 l0bl14 vdd x644 x644b CELLD r1=900e3 r0=10000e3
xl0b14c645 l0bl14 vdd x645 x645b CELLD r1=10000e3 r0=900e3
xl0b14c646 l0bl14 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b14c647 l0bl14 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b14c648 l0bl14 vdd x648 x648b CELLD r1=10000e3 r0=900e3
xl0b14c649 l0bl14 vdd x649 x649b CELLD r1=900e3 r0=10000e3
xl0b14c650 l0bl14 vdd x650 x650b CELLD r1=900e3 r0=10000e3
xl0b14c651 l0bl14 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b14c652 l0bl14 vdd x652 x652b CELLD r1=900e3 r0=10000e3
xl0b14c653 l0bl14 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b14c654 l0bl14 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b14c655 l0bl14 vdd x655 x655b CELLD r1=900e3 r0=10000e3
xl0b14c656 l0bl14 vdd x656 x656b CELLD r1=900e3 r0=10000e3
xl0b14c657 l0bl14 vdd x657 x657b CELLD r1=900e3 r0=10000e3
xl0b14c658 l0bl14 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b14c659 l0bl14 vdd x659 x659b CELLD r1=900e3 r0=10000e3
xl0b14c660 l0bl14 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b14c661 l0bl14 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b14c662 l0bl14 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b14c663 l0bl14 vdd x663 x663b CELLD r1=10000e3 r0=900e3
xl0b14c664 l0bl14 vdd x664 x664b CELLD r1=10000e3 r0=900e3
xl0b14c665 l0bl14 vdd x665 x665b CELLD r1=10000e3 r0=900e3
xl0b14c666 l0bl14 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b14c667 l0bl14 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b14c668 l0bl14 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b14c669 l0bl14 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b14c670 l0bl14 vdd x670 x670b CELLD r1=10000e3 r0=900e3
xl0b14c671 l0bl14 vdd x671 x671b CELLD r1=10000e3 r0=900e3
xl0b14c672 l0bl14 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b14c673 l0bl14 vdd x673 x673b CELLD r1=10000e3 r0=900e3
xl0b14c674 l0bl14 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b14c675 l0bl14 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b14c676 l0bl14 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b14c677 l0bl14 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b14c678 l0bl14 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b14c679 l0bl14 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b14c680 l0bl14 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b14c681 l0bl14 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b14c682 l0bl14 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b14c683 l0bl14 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b14c684 l0bl14 vdd x684 x684b CELLD r1=900e3 r0=10000e3
xl0b14c685 l0bl14 vdd x685 x685b CELLD r1=900e3 r0=10000e3
xl0b14c686 l0bl14 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b14c687 l0bl14 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b14c688 l0bl14 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b14c689 l0bl14 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b14c690 l0bl14 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b14c691 l0bl14 vdd x691 x691b CELLD r1=10000e3 r0=900e3
xl0b14c692 l0bl14 vdd x692 x692b CELLD r1=10000e3 r0=900e3
xl0b14c693 l0bl14 vdd x693 x693b CELLD r1=10000e3 r0=900e3
xl0b14c694 l0bl14 vdd x694 x694b CELLD r1=10000e3 r0=900e3
xl0b14c695 l0bl14 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b14c696 l0bl14 vdd x696 x696b CELLD r1=10000e3 r0=900e3
xl0b14c697 l0bl14 vdd x697 x697b CELLD r1=10000e3 r0=900e3
xl0b14c698 l0bl14 vdd x698 x698b CELLD r1=10000e3 r0=900e3
xl0b14c699 l0bl14 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b14c700 l0bl14 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b14c701 l0bl14 vdd x701 x701b CELLD r1=10000e3 r0=900e3
xl0b14c702 l0bl14 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b14c703 l0bl14 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b14c704 l0bl14 vdd x704 x704b CELLD r1=10000e3 r0=900e3
xl0b14c705 l0bl14 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b14c706 l0bl14 vdd x706 x706b CELLD r1=10000e3 r0=900e3
xl0b14c707 l0bl14 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b14c708 l0bl14 vdd x708 x708b CELLD r1=10000e3 r0=900e3
xl0b14c709 l0bl14 vdd x709 x709b CELLD r1=10000e3 r0=900e3
xl0b14c710 l0bl14 vdd x710 x710b CELLD r1=10000e3 r0=900e3
xl0b14c711 l0bl14 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b14c712 l0bl14 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b14c713 l0bl14 vdd x713 x713b CELLD r1=10000e3 r0=900e3
xl0b14c714 l0bl14 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b14c715 l0bl14 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b14c716 l0bl14 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b14c717 l0bl14 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b14c718 l0bl14 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b14c719 l0bl14 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b14c720 l0bl14 vdd x720 x720b CELLD r1=10000e3 r0=900e3
xl0b14c721 l0bl14 vdd x721 x721b CELLD r1=10000e3 r0=900e3
xl0b14c722 l0bl14 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b14c723 l0bl14 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b14c724 l0bl14 vdd x724 x724b CELLD r1=10000e3 r0=900e3
xl0b14c725 l0bl14 vdd x725 x725b CELLD r1=10000e3 r0=900e3
xl0b14c726 l0bl14 vdd x726 x726b CELLD r1=10000e3 r0=900e3
xl0b14c727 l0bl14 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b14c728 l0bl14 vdd x728 x728b CELLD r1=10000e3 r0=900e3
xl0b14c729 l0bl14 vdd x729 x729b CELLD r1=10000e3 r0=900e3
xl0b14c730 l0bl14 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b14c731 l0bl14 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b14c732 l0bl14 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b14c733 l0bl14 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b14c734 l0bl14 vdd x734 x734b CELLD r1=10000e3 r0=900e3
xl0b14c735 l0bl14 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b14c736 l0bl14 vdd x736 x736b CELLD r1=10000e3 r0=900e3
xl0b14c737 l0bl14 vdd x737 x737b CELLD r1=10000e3 r0=900e3
xl0b14c738 l0bl14 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b14c739 l0bl14 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b14c740 l0bl14 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b14c741 l0bl14 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b14c742 l0bl14 vdd x742 x742b CELLD r1=10000e3 r0=900e3
xl0b14c743 l0bl14 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b14c744 l0bl14 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b14c745 l0bl14 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b14c746 l0bl14 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b14c747 l0bl14 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b14c748 l0bl14 vdd x748 x748b CELLD r1=10000e3 r0=900e3
xl0b14c749 l0bl14 vdd x749 x749b CELLD r1=10000e3 r0=900e3
xl0b14c750 l0bl14 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b14c751 l0bl14 vdd x751 x751b CELLD r1=10000e3 r0=900e3
xl0b14c752 l0bl14 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b14c753 l0bl14 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b14c754 l0bl14 vdd x754 x754b CELLD r1=10000e3 r0=900e3
xl0b14c755 l0bl14 vdd x755 x755b CELLD r1=10000e3 r0=900e3
xl0b14c756 l0bl14 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b14c757 l0bl14 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b14c758 l0bl14 vdd x758 x758b CELLD r1=10000e3 r0=900e3
xl0b14c759 l0bl14 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b14c760 l0bl14 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b14c761 l0bl14 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b14c762 l0bl14 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b14c763 l0bl14 vdd x763 x763b CELLD r1=10000e3 r0=900e3
xl0b14c764 l0bl14 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b14c765 l0bl14 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b14c766 l0bl14 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b14c767 l0bl14 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b14c768 l0bl14 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b14c769 l0bl14 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b14c770 l0bl14 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b14c771 l0bl14 vdd x771 x771b CELLD r1=10000e3 r0=900e3
xl0b14c772 l0bl14 vdd x772 x772b CELLD r1=10000e3 r0=900e3
xl0b14c773 l0bl14 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b14c774 l0bl14 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b14c775 l0bl14 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b14c776 l0bl14 vdd x776 x776b CELLD r1=10000e3 r0=900e3
xl0b14c777 l0bl14 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b14c778 l0bl14 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b14c779 l0bl14 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b14c780 l0bl14 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b14c781 l0bl14 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b14c782 l0bl14 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b14c783 l0bl14 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b15c0 l0bl15 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b15c1 l0bl15 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b15c2 l0bl15 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b15c3 l0bl15 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b15c4 l0bl15 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b15c5 l0bl15 vdd x5 x5b CELLD r1=10000e3 r0=900e3
xl0b15c6 l0bl15 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b15c7 l0bl15 vdd x7 x7b CELLD r1=900e3 r0=10000e3
xl0b15c8 l0bl15 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b15c9 l0bl15 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b15c10 l0bl15 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b15c11 l0bl15 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b15c12 l0bl15 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b15c13 l0bl15 vdd x13 x13b CELLD r1=10000e3 r0=900e3
xl0b15c14 l0bl15 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b15c15 l0bl15 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b15c16 l0bl15 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b15c17 l0bl15 vdd x17 x17b CELLD r1=10000e3 r0=900e3
xl0b15c18 l0bl15 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b15c19 l0bl15 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b15c20 l0bl15 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b15c21 l0bl15 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b15c22 l0bl15 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b15c23 l0bl15 vdd x23 x23b CELLD r1=10000e3 r0=900e3
xl0b15c24 l0bl15 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b15c25 l0bl15 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b15c26 l0bl15 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b15c27 l0bl15 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b15c28 l0bl15 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b15c29 l0bl15 vdd x29 x29b CELLD r1=10000e3 r0=900e3
xl0b15c30 l0bl15 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b15c31 l0bl15 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b15c32 l0bl15 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b15c33 l0bl15 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b15c34 l0bl15 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b15c35 l0bl15 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b15c36 l0bl15 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b15c37 l0bl15 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b15c38 l0bl15 vdd x38 x38b CELLD r1=10000e3 r0=900e3
xl0b15c39 l0bl15 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b15c40 l0bl15 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b15c41 l0bl15 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b15c42 l0bl15 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b15c43 l0bl15 vdd x43 x43b CELLD r1=10000e3 r0=900e3
xl0b15c44 l0bl15 vdd x44 x44b CELLD r1=10000e3 r0=900e3
xl0b15c45 l0bl15 vdd x45 x45b CELLD r1=900e3 r0=10000e3
xl0b15c46 l0bl15 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b15c47 l0bl15 vdd x47 x47b CELLD r1=900e3 r0=10000e3
xl0b15c48 l0bl15 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b15c49 l0bl15 vdd x49 x49b CELLD r1=900e3 r0=10000e3
xl0b15c50 l0bl15 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b15c51 l0bl15 vdd x51 x51b CELLD r1=900e3 r0=10000e3
xl0b15c52 l0bl15 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b15c53 l0bl15 vdd x53 x53b CELLD r1=900e3 r0=10000e3
xl0b15c54 l0bl15 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b15c55 l0bl15 vdd x55 x55b CELLD r1=900e3 r0=10000e3
xl0b15c56 l0bl15 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b15c57 l0bl15 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b15c58 l0bl15 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b15c59 l0bl15 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b15c60 l0bl15 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b15c61 l0bl15 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b15c62 l0bl15 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b15c63 l0bl15 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b15c64 l0bl15 vdd x64 x64b CELLD r1=900e3 r0=10000e3
xl0b15c65 l0bl15 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b15c66 l0bl15 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b15c67 l0bl15 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b15c68 l0bl15 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b15c69 l0bl15 vdd x69 x69b CELLD r1=900e3 r0=10000e3
xl0b15c70 l0bl15 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b15c71 l0bl15 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b15c72 l0bl15 vdd x72 x72b CELLD r1=900e3 r0=10000e3
xl0b15c73 l0bl15 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b15c74 l0bl15 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b15c75 l0bl15 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b15c76 l0bl15 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b15c77 l0bl15 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b15c78 l0bl15 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b15c79 l0bl15 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b15c80 l0bl15 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b15c81 l0bl15 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b15c82 l0bl15 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b15c83 l0bl15 vdd x83 x83b CELLD r1=900e3 r0=10000e3
xl0b15c84 l0bl15 vdd x84 x84b CELLD r1=900e3 r0=10000e3
xl0b15c85 l0bl15 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b15c86 l0bl15 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b15c87 l0bl15 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b15c88 l0bl15 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b15c89 l0bl15 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b15c90 l0bl15 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b15c91 l0bl15 vdd x91 x91b CELLD r1=900e3 r0=10000e3
xl0b15c92 l0bl15 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b15c93 l0bl15 vdd x93 x93b CELLD r1=900e3 r0=10000e3
xl0b15c94 l0bl15 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b15c95 l0bl15 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b15c96 l0bl15 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b15c97 l0bl15 vdd x97 x97b CELLD r1=900e3 r0=10000e3
xl0b15c98 l0bl15 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b15c99 l0bl15 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b15c100 l0bl15 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b15c101 l0bl15 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b15c102 l0bl15 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b15c103 l0bl15 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b15c104 l0bl15 vdd x104 x104b CELLD r1=900e3 r0=10000e3
xl0b15c105 l0bl15 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b15c106 l0bl15 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b15c107 l0bl15 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b15c108 l0bl15 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b15c109 l0bl15 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b15c110 l0bl15 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b15c111 l0bl15 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b15c112 l0bl15 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b15c113 l0bl15 vdd x113 x113b CELLD r1=900e3 r0=10000e3
xl0b15c114 l0bl15 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b15c115 l0bl15 vdd x115 x115b CELLD r1=900e3 r0=10000e3
xl0b15c116 l0bl15 vdd x116 x116b CELLD r1=10000e3 r0=900e3
xl0b15c117 l0bl15 vdd x117 x117b CELLD r1=900e3 r0=10000e3
xl0b15c118 l0bl15 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b15c119 l0bl15 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b15c120 l0bl15 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b15c121 l0bl15 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b15c122 l0bl15 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b15c123 l0bl15 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b15c124 l0bl15 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b15c125 l0bl15 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b15c126 l0bl15 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b15c127 l0bl15 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b15c128 l0bl15 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b15c129 l0bl15 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b15c130 l0bl15 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b15c131 l0bl15 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b15c132 l0bl15 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b15c133 l0bl15 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b15c134 l0bl15 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b15c135 l0bl15 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b15c136 l0bl15 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b15c137 l0bl15 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b15c138 l0bl15 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b15c139 l0bl15 vdd x139 x139b CELLD r1=900e3 r0=10000e3
xl0b15c140 l0bl15 vdd x140 x140b CELLD r1=900e3 r0=10000e3
xl0b15c141 l0bl15 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b15c142 l0bl15 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b15c143 l0bl15 vdd x143 x143b CELLD r1=10000e3 r0=900e3
xl0b15c144 l0bl15 vdd x144 x144b CELLD r1=900e3 r0=10000e3
xl0b15c145 l0bl15 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b15c146 l0bl15 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b15c147 l0bl15 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b15c148 l0bl15 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b15c149 l0bl15 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b15c150 l0bl15 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b15c151 l0bl15 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b15c152 l0bl15 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b15c153 l0bl15 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b15c154 l0bl15 vdd x154 x154b CELLD r1=10000e3 r0=900e3
xl0b15c155 l0bl15 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b15c156 l0bl15 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b15c157 l0bl15 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b15c158 l0bl15 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b15c159 l0bl15 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b15c160 l0bl15 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b15c161 l0bl15 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b15c162 l0bl15 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b15c163 l0bl15 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b15c164 l0bl15 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b15c165 l0bl15 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b15c166 l0bl15 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b15c167 l0bl15 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b15c168 l0bl15 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b15c169 l0bl15 vdd x169 x169b CELLD r1=10000e3 r0=900e3
xl0b15c170 l0bl15 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b15c171 l0bl15 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b15c172 l0bl15 vdd x172 x172b CELLD r1=10000e3 r0=900e3
xl0b15c173 l0bl15 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b15c174 l0bl15 vdd x174 x174b CELLD r1=10000e3 r0=900e3
xl0b15c175 l0bl15 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b15c176 l0bl15 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b15c177 l0bl15 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b15c178 l0bl15 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b15c179 l0bl15 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b15c180 l0bl15 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b15c181 l0bl15 vdd x181 x181b CELLD r1=10000e3 r0=900e3
xl0b15c182 l0bl15 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b15c183 l0bl15 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b15c184 l0bl15 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b15c185 l0bl15 vdd x185 x185b CELLD r1=10000e3 r0=900e3
xl0b15c186 l0bl15 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b15c187 l0bl15 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b15c188 l0bl15 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b15c189 l0bl15 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b15c190 l0bl15 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b15c191 l0bl15 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b15c192 l0bl15 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b15c193 l0bl15 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b15c194 l0bl15 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b15c195 l0bl15 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b15c196 l0bl15 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b15c197 l0bl15 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b15c198 l0bl15 vdd x198 x198b CELLD r1=900e3 r0=10000e3
xl0b15c199 l0bl15 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b15c200 l0bl15 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b15c201 l0bl15 vdd x201 x201b CELLD r1=10000e3 r0=900e3
xl0b15c202 l0bl15 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b15c203 l0bl15 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b15c204 l0bl15 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b15c205 l0bl15 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b15c206 l0bl15 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b15c207 l0bl15 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b15c208 l0bl15 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b15c209 l0bl15 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b15c210 l0bl15 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b15c211 l0bl15 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b15c212 l0bl15 vdd x212 x212b CELLD r1=10000e3 r0=900e3
xl0b15c213 l0bl15 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b15c214 l0bl15 vdd x214 x214b CELLD r1=10000e3 r0=900e3
xl0b15c215 l0bl15 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b15c216 l0bl15 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b15c217 l0bl15 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b15c218 l0bl15 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b15c219 l0bl15 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b15c220 l0bl15 vdd x220 x220b CELLD r1=900e3 r0=10000e3
xl0b15c221 l0bl15 vdd x221 x221b CELLD r1=900e3 r0=10000e3
xl0b15c222 l0bl15 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b15c223 l0bl15 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b15c224 l0bl15 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b15c225 l0bl15 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b15c226 l0bl15 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b15c227 l0bl15 vdd x227 x227b CELLD r1=10000e3 r0=900e3
xl0b15c228 l0bl15 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b15c229 l0bl15 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b15c230 l0bl15 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b15c231 l0bl15 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b15c232 l0bl15 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b15c233 l0bl15 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b15c234 l0bl15 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b15c235 l0bl15 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b15c236 l0bl15 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b15c237 l0bl15 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b15c238 l0bl15 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b15c239 l0bl15 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b15c240 l0bl15 vdd x240 x240b CELLD r1=10000e3 r0=900e3
xl0b15c241 l0bl15 vdd x241 x241b CELLD r1=10000e3 r0=900e3
xl0b15c242 l0bl15 vdd x242 x242b CELLD r1=10000e3 r0=900e3
xl0b15c243 l0bl15 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b15c244 l0bl15 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b15c245 l0bl15 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b15c246 l0bl15 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b15c247 l0bl15 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b15c248 l0bl15 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b15c249 l0bl15 vdd x249 x249b CELLD r1=900e3 r0=10000e3
xl0b15c250 l0bl15 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b15c251 l0bl15 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b15c252 l0bl15 vdd x252 x252b CELLD r1=900e3 r0=10000e3
xl0b15c253 l0bl15 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b15c254 l0bl15 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b15c255 l0bl15 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b15c256 l0bl15 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b15c257 l0bl15 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b15c258 l0bl15 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b15c259 l0bl15 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b15c260 l0bl15 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b15c261 l0bl15 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b15c262 l0bl15 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b15c263 l0bl15 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b15c264 l0bl15 vdd x264 x264b CELLD r1=10000e3 r0=900e3
xl0b15c265 l0bl15 vdd x265 x265b CELLD r1=10000e3 r0=900e3
xl0b15c266 l0bl15 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b15c267 l0bl15 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b15c268 l0bl15 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b15c269 l0bl15 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b15c270 l0bl15 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b15c271 l0bl15 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b15c272 l0bl15 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b15c273 l0bl15 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b15c274 l0bl15 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b15c275 l0bl15 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b15c276 l0bl15 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b15c277 l0bl15 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b15c278 l0bl15 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b15c279 l0bl15 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b15c280 l0bl15 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b15c281 l0bl15 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b15c282 l0bl15 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b15c283 l0bl15 vdd x283 x283b CELLD r1=10000e3 r0=900e3
xl0b15c284 l0bl15 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b15c285 l0bl15 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b15c286 l0bl15 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b15c287 l0bl15 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b15c288 l0bl15 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b15c289 l0bl15 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b15c290 l0bl15 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b15c291 l0bl15 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b15c292 l0bl15 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b15c293 l0bl15 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b15c294 l0bl15 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b15c295 l0bl15 vdd x295 x295b CELLD r1=10000e3 r0=900e3
xl0b15c296 l0bl15 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b15c297 l0bl15 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b15c298 l0bl15 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b15c299 l0bl15 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b15c300 l0bl15 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b15c301 l0bl15 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b15c302 l0bl15 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b15c303 l0bl15 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b15c304 l0bl15 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b15c305 l0bl15 vdd x305 x305b CELLD r1=900e3 r0=10000e3
xl0b15c306 l0bl15 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b15c307 l0bl15 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b15c308 l0bl15 vdd x308 x308b CELLD r1=10000e3 r0=900e3
xl0b15c309 l0bl15 vdd x309 x309b CELLD r1=10000e3 r0=900e3
xl0b15c310 l0bl15 vdd x310 x310b CELLD r1=900e3 r0=10000e3
xl0b15c311 l0bl15 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b15c312 l0bl15 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b15c313 l0bl15 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b15c314 l0bl15 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b15c315 l0bl15 vdd x315 x315b CELLD r1=900e3 r0=10000e3
xl0b15c316 l0bl15 vdd x316 x316b CELLD r1=900e3 r0=10000e3
xl0b15c317 l0bl15 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b15c318 l0bl15 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b15c319 l0bl15 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b15c320 l0bl15 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b15c321 l0bl15 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b15c322 l0bl15 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b15c323 l0bl15 vdd x323 x323b CELLD r1=10000e3 r0=900e3
xl0b15c324 l0bl15 vdd x324 x324b CELLD r1=10000e3 r0=900e3
xl0b15c325 l0bl15 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b15c326 l0bl15 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b15c327 l0bl15 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b15c328 l0bl15 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b15c329 l0bl15 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b15c330 l0bl15 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b15c331 l0bl15 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b15c332 l0bl15 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b15c333 l0bl15 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b15c334 l0bl15 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b15c335 l0bl15 vdd x335 x335b CELLD r1=10000e3 r0=900e3
xl0b15c336 l0bl15 vdd x336 x336b CELLD r1=900e3 r0=10000e3
xl0b15c337 l0bl15 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b15c338 l0bl15 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b15c339 l0bl15 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b15c340 l0bl15 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b15c341 l0bl15 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b15c342 l0bl15 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b15c343 l0bl15 vdd x343 x343b CELLD r1=900e3 r0=10000e3
xl0b15c344 l0bl15 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b15c345 l0bl15 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b15c346 l0bl15 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b15c347 l0bl15 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b15c348 l0bl15 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b15c349 l0bl15 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b15c350 l0bl15 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b15c351 l0bl15 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b15c352 l0bl15 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b15c353 l0bl15 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b15c354 l0bl15 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b15c355 l0bl15 vdd x355 x355b CELLD r1=900e3 r0=10000e3
xl0b15c356 l0bl15 vdd x356 x356b CELLD r1=900e3 r0=10000e3
xl0b15c357 l0bl15 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b15c358 l0bl15 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b15c359 l0bl15 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b15c360 l0bl15 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b15c361 l0bl15 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b15c362 l0bl15 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b15c363 l0bl15 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b15c364 l0bl15 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b15c365 l0bl15 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b15c366 l0bl15 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b15c367 l0bl15 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b15c368 l0bl15 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b15c369 l0bl15 vdd x369 x369b CELLD r1=900e3 r0=10000e3
xl0b15c370 l0bl15 vdd x370 x370b CELLD r1=900e3 r0=10000e3
xl0b15c371 l0bl15 vdd x371 x371b CELLD r1=900e3 r0=10000e3
xl0b15c372 l0bl15 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b15c373 l0bl15 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b15c374 l0bl15 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b15c375 l0bl15 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b15c376 l0bl15 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b15c377 l0bl15 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b15c378 l0bl15 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b15c379 l0bl15 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b15c380 l0bl15 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b15c381 l0bl15 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b15c382 l0bl15 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b15c383 l0bl15 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b15c384 l0bl15 vdd x384 x384b CELLD r1=900e3 r0=10000e3
xl0b15c385 l0bl15 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b15c386 l0bl15 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b15c387 l0bl15 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b15c388 l0bl15 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b15c389 l0bl15 vdd x389 x389b CELLD r1=10000e3 r0=900e3
xl0b15c390 l0bl15 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b15c391 l0bl15 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b15c392 l0bl15 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b15c393 l0bl15 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b15c394 l0bl15 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b15c395 l0bl15 vdd x395 x395b CELLD r1=900e3 r0=10000e3
xl0b15c396 l0bl15 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b15c397 l0bl15 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b15c398 l0bl15 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b15c399 l0bl15 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b15c400 l0bl15 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b15c401 l0bl15 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b15c402 l0bl15 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b15c403 l0bl15 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b15c404 l0bl15 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b15c405 l0bl15 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b15c406 l0bl15 vdd x406 x406b CELLD r1=10000e3 r0=900e3
xl0b15c407 l0bl15 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b15c408 l0bl15 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b15c409 l0bl15 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b15c410 l0bl15 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b15c411 l0bl15 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b15c412 l0bl15 vdd x412 x412b CELLD r1=900e3 r0=10000e3
xl0b15c413 l0bl15 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b15c414 l0bl15 vdd x414 x414b CELLD r1=900e3 r0=10000e3
xl0b15c415 l0bl15 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b15c416 l0bl15 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b15c417 l0bl15 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b15c418 l0bl15 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b15c419 l0bl15 vdd x419 x419b CELLD r1=900e3 r0=10000e3
xl0b15c420 l0bl15 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b15c421 l0bl15 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b15c422 l0bl15 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b15c423 l0bl15 vdd x423 x423b CELLD r1=900e3 r0=10000e3
xl0b15c424 l0bl15 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b15c425 l0bl15 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b15c426 l0bl15 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b15c427 l0bl15 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b15c428 l0bl15 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b15c429 l0bl15 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b15c430 l0bl15 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b15c431 l0bl15 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b15c432 l0bl15 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b15c433 l0bl15 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b15c434 l0bl15 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b15c435 l0bl15 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b15c436 l0bl15 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b15c437 l0bl15 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b15c438 l0bl15 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b15c439 l0bl15 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b15c440 l0bl15 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b15c441 l0bl15 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b15c442 l0bl15 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b15c443 l0bl15 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b15c444 l0bl15 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b15c445 l0bl15 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b15c446 l0bl15 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b15c447 l0bl15 vdd x447 x447b CELLD r1=10000e3 r0=900e3
xl0b15c448 l0bl15 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b15c449 l0bl15 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b15c450 l0bl15 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b15c451 l0bl15 vdd x451 x451b CELLD r1=900e3 r0=10000e3
xl0b15c452 l0bl15 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b15c453 l0bl15 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b15c454 l0bl15 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b15c455 l0bl15 vdd x455 x455b CELLD r1=900e3 r0=10000e3
xl0b15c456 l0bl15 vdd x456 x456b CELLD r1=900e3 r0=10000e3
xl0b15c457 l0bl15 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b15c458 l0bl15 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b15c459 l0bl15 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b15c460 l0bl15 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b15c461 l0bl15 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b15c462 l0bl15 vdd x462 x462b CELLD r1=10000e3 r0=900e3
xl0b15c463 l0bl15 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b15c464 l0bl15 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b15c465 l0bl15 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b15c466 l0bl15 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b15c467 l0bl15 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b15c468 l0bl15 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b15c469 l0bl15 vdd x469 x469b CELLD r1=900e3 r0=10000e3
xl0b15c470 l0bl15 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b15c471 l0bl15 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b15c472 l0bl15 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b15c473 l0bl15 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b15c474 l0bl15 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b15c475 l0bl15 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b15c476 l0bl15 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b15c477 l0bl15 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b15c478 l0bl15 vdd x478 x478b CELLD r1=900e3 r0=10000e3
xl0b15c479 l0bl15 vdd x479 x479b CELLD r1=900e3 r0=10000e3
xl0b15c480 l0bl15 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b15c481 l0bl15 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b15c482 l0bl15 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b15c483 l0bl15 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b15c484 l0bl15 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b15c485 l0bl15 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b15c486 l0bl15 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b15c487 l0bl15 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b15c488 l0bl15 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b15c489 l0bl15 vdd x489 x489b CELLD r1=10000e3 r0=900e3
xl0b15c490 l0bl15 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b15c491 l0bl15 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b15c492 l0bl15 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b15c493 l0bl15 vdd x493 x493b CELLD r1=10000e3 r0=900e3
xl0b15c494 l0bl15 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b15c495 l0bl15 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b15c496 l0bl15 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b15c497 l0bl15 vdd x497 x497b CELLD r1=900e3 r0=10000e3
xl0b15c498 l0bl15 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b15c499 l0bl15 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b15c500 l0bl15 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b15c501 l0bl15 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b15c502 l0bl15 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b15c503 l0bl15 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b15c504 l0bl15 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b15c505 l0bl15 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b15c506 l0bl15 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b15c507 l0bl15 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b15c508 l0bl15 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b15c509 l0bl15 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b15c510 l0bl15 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b15c511 l0bl15 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b15c512 l0bl15 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b15c513 l0bl15 vdd x513 x513b CELLD r1=10000e3 r0=900e3
xl0b15c514 l0bl15 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b15c515 l0bl15 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b15c516 l0bl15 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b15c517 l0bl15 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b15c518 l0bl15 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b15c519 l0bl15 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b15c520 l0bl15 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b15c521 l0bl15 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b15c522 l0bl15 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b15c523 l0bl15 vdd x523 x523b CELLD r1=900e3 r0=10000e3
xl0b15c524 l0bl15 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b15c525 l0bl15 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b15c526 l0bl15 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b15c527 l0bl15 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b15c528 l0bl15 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b15c529 l0bl15 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b15c530 l0bl15 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b15c531 l0bl15 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b15c532 l0bl15 vdd x532 x532b CELLD r1=10000e3 r0=900e3
xl0b15c533 l0bl15 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b15c534 l0bl15 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b15c535 l0bl15 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b15c536 l0bl15 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b15c537 l0bl15 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b15c538 l0bl15 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b15c539 l0bl15 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b15c540 l0bl15 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b15c541 l0bl15 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b15c542 l0bl15 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b15c543 l0bl15 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b15c544 l0bl15 vdd x544 x544b CELLD r1=10000e3 r0=900e3
xl0b15c545 l0bl15 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b15c546 l0bl15 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b15c547 l0bl15 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b15c548 l0bl15 vdd x548 x548b CELLD r1=900e3 r0=10000e3
xl0b15c549 l0bl15 vdd x549 x549b CELLD r1=900e3 r0=10000e3
xl0b15c550 l0bl15 vdd x550 x550b CELLD r1=900e3 r0=10000e3
xl0b15c551 l0bl15 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b15c552 l0bl15 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b15c553 l0bl15 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b15c554 l0bl15 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b15c555 l0bl15 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b15c556 l0bl15 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b15c557 l0bl15 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b15c558 l0bl15 vdd x558 x558b CELLD r1=10000e3 r0=900e3
xl0b15c559 l0bl15 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b15c560 l0bl15 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b15c561 l0bl15 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b15c562 l0bl15 vdd x562 x562b CELLD r1=900e3 r0=10000e3
xl0b15c563 l0bl15 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b15c564 l0bl15 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b15c565 l0bl15 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b15c566 l0bl15 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b15c567 l0bl15 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b15c568 l0bl15 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b15c569 l0bl15 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b15c570 l0bl15 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b15c571 l0bl15 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b15c572 l0bl15 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b15c573 l0bl15 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b15c574 l0bl15 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b15c575 l0bl15 vdd x575 x575b CELLD r1=900e3 r0=10000e3
xl0b15c576 l0bl15 vdd x576 x576b CELLD r1=900e3 r0=10000e3
xl0b15c577 l0bl15 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b15c578 l0bl15 vdd x578 x578b CELLD r1=900e3 r0=10000e3
xl0b15c579 l0bl15 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b15c580 l0bl15 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b15c581 l0bl15 vdd x581 x581b CELLD r1=10000e3 r0=900e3
xl0b15c582 l0bl15 vdd x582 x582b CELLD r1=10000e3 r0=900e3
xl0b15c583 l0bl15 vdd x583 x583b CELLD r1=10000e3 r0=900e3
xl0b15c584 l0bl15 vdd x584 x584b CELLD r1=10000e3 r0=900e3
xl0b15c585 l0bl15 vdd x585 x585b CELLD r1=10000e3 r0=900e3
xl0b15c586 l0bl15 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b15c587 l0bl15 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b15c588 l0bl15 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b15c589 l0bl15 vdd x589 x589b CELLD r1=10000e3 r0=900e3
xl0b15c590 l0bl15 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b15c591 l0bl15 vdd x591 x591b CELLD r1=900e3 r0=10000e3
xl0b15c592 l0bl15 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b15c593 l0bl15 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b15c594 l0bl15 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b15c595 l0bl15 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b15c596 l0bl15 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b15c597 l0bl15 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b15c598 l0bl15 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b15c599 l0bl15 vdd x599 x599b CELLD r1=900e3 r0=10000e3
xl0b15c600 l0bl15 vdd x600 x600b CELLD r1=900e3 r0=10000e3
xl0b15c601 l0bl15 vdd x601 x601b CELLD r1=900e3 r0=10000e3
xl0b15c602 l0bl15 vdd x602 x602b CELLD r1=900e3 r0=10000e3
xl0b15c603 l0bl15 vdd x603 x603b CELLD r1=900e3 r0=10000e3
xl0b15c604 l0bl15 vdd x604 x604b CELLD r1=900e3 r0=10000e3
xl0b15c605 l0bl15 vdd x605 x605b CELLD r1=900e3 r0=10000e3
xl0b15c606 l0bl15 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b15c607 l0bl15 vdd x607 x607b CELLD r1=10000e3 r0=900e3
xl0b15c608 l0bl15 vdd x608 x608b CELLD r1=10000e3 r0=900e3
xl0b15c609 l0bl15 vdd x609 x609b CELLD r1=10000e3 r0=900e3
xl0b15c610 l0bl15 vdd x610 x610b CELLD r1=10000e3 r0=900e3
xl0b15c611 l0bl15 vdd x611 x611b CELLD r1=10000e3 r0=900e3
xl0b15c612 l0bl15 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b15c613 l0bl15 vdd x613 x613b CELLD r1=900e3 r0=10000e3
xl0b15c614 l0bl15 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b15c615 l0bl15 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b15c616 l0bl15 vdd x616 x616b CELLD r1=10000e3 r0=900e3
xl0b15c617 l0bl15 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b15c618 l0bl15 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b15c619 l0bl15 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b15c620 l0bl15 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b15c621 l0bl15 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b15c622 l0bl15 vdd x622 x622b CELLD r1=10000e3 r0=900e3
xl0b15c623 l0bl15 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b15c624 l0bl15 vdd x624 x624b CELLD r1=10000e3 r0=900e3
xl0b15c625 l0bl15 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b15c626 l0bl15 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b15c627 l0bl15 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b15c628 l0bl15 vdd x628 x628b CELLD r1=900e3 r0=10000e3
xl0b15c629 l0bl15 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b15c630 l0bl15 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b15c631 l0bl15 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b15c632 l0bl15 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b15c633 l0bl15 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b15c634 l0bl15 vdd x634 x634b CELLD r1=10000e3 r0=900e3
xl0b15c635 l0bl15 vdd x635 x635b CELLD r1=10000e3 r0=900e3
xl0b15c636 l0bl15 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b15c637 l0bl15 vdd x637 x637b CELLD r1=10000e3 r0=900e3
xl0b15c638 l0bl15 vdd x638 x638b CELLD r1=10000e3 r0=900e3
xl0b15c639 l0bl15 vdd x639 x639b CELLD r1=10000e3 r0=900e3
xl0b15c640 l0bl15 vdd x640 x640b CELLD r1=10000e3 r0=900e3
xl0b15c641 l0bl15 vdd x641 x641b CELLD r1=10000e3 r0=900e3
xl0b15c642 l0bl15 vdd x642 x642b CELLD r1=10000e3 r0=900e3
xl0b15c643 l0bl15 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b15c644 l0bl15 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b15c645 l0bl15 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b15c646 l0bl15 vdd x646 x646b CELLD r1=900e3 r0=10000e3
xl0b15c647 l0bl15 vdd x647 x647b CELLD r1=900e3 r0=10000e3
xl0b15c648 l0bl15 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b15c649 l0bl15 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b15c650 l0bl15 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b15c651 l0bl15 vdd x651 x651b CELLD r1=10000e3 r0=900e3
xl0b15c652 l0bl15 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b15c653 l0bl15 vdd x653 x653b CELLD r1=10000e3 r0=900e3
xl0b15c654 l0bl15 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b15c655 l0bl15 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b15c656 l0bl15 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b15c657 l0bl15 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b15c658 l0bl15 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b15c659 l0bl15 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b15c660 l0bl15 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b15c661 l0bl15 vdd x661 x661b CELLD r1=10000e3 r0=900e3
xl0b15c662 l0bl15 vdd x662 x662b CELLD r1=10000e3 r0=900e3
xl0b15c663 l0bl15 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b15c664 l0bl15 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b15c665 l0bl15 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b15c666 l0bl15 vdd x666 x666b CELLD r1=900e3 r0=10000e3
xl0b15c667 l0bl15 vdd x667 x667b CELLD r1=900e3 r0=10000e3
xl0b15c668 l0bl15 vdd x668 x668b CELLD r1=10000e3 r0=900e3
xl0b15c669 l0bl15 vdd x669 x669b CELLD r1=10000e3 r0=900e3
xl0b15c670 l0bl15 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b15c671 l0bl15 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b15c672 l0bl15 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b15c673 l0bl15 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b15c674 l0bl15 vdd x674 x674b CELLD r1=900e3 r0=10000e3
xl0b15c675 l0bl15 vdd x675 x675b CELLD r1=900e3 r0=10000e3
xl0b15c676 l0bl15 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b15c677 l0bl15 vdd x677 x677b CELLD r1=10000e3 r0=900e3
xl0b15c678 l0bl15 vdd x678 x678b CELLD r1=10000e3 r0=900e3
xl0b15c679 l0bl15 vdd x679 x679b CELLD r1=10000e3 r0=900e3
xl0b15c680 l0bl15 vdd x680 x680b CELLD r1=10000e3 r0=900e3
xl0b15c681 l0bl15 vdd x681 x681b CELLD r1=10000e3 r0=900e3
xl0b15c682 l0bl15 vdd x682 x682b CELLD r1=10000e3 r0=900e3
xl0b15c683 l0bl15 vdd x683 x683b CELLD r1=900e3 r0=10000e3
xl0b15c684 l0bl15 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b15c685 l0bl15 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b15c686 l0bl15 vdd x686 x686b CELLD r1=10000e3 r0=900e3
xl0b15c687 l0bl15 vdd x687 x687b CELLD r1=10000e3 r0=900e3
xl0b15c688 l0bl15 vdd x688 x688b CELLD r1=10000e3 r0=900e3
xl0b15c689 l0bl15 vdd x689 x689b CELLD r1=10000e3 r0=900e3
xl0b15c690 l0bl15 vdd x690 x690b CELLD r1=10000e3 r0=900e3
xl0b15c691 l0bl15 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b15c692 l0bl15 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b15c693 l0bl15 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b15c694 l0bl15 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b15c695 l0bl15 vdd x695 x695b CELLD r1=10000e3 r0=900e3
xl0b15c696 l0bl15 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b15c697 l0bl15 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b15c698 l0bl15 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b15c699 l0bl15 vdd x699 x699b CELLD r1=900e3 r0=10000e3
xl0b15c700 l0bl15 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b15c701 l0bl15 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b15c702 l0bl15 vdd x702 x702b CELLD r1=900e3 r0=10000e3
xl0b15c703 l0bl15 vdd x703 x703b CELLD r1=10000e3 r0=900e3
xl0b15c704 l0bl15 vdd x704 x704b CELLD r1=900e3 r0=10000e3
xl0b15c705 l0bl15 vdd x705 x705b CELLD r1=10000e3 r0=900e3
xl0b15c706 l0bl15 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b15c707 l0bl15 vdd x707 x707b CELLD r1=10000e3 r0=900e3
xl0b15c708 l0bl15 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b15c709 l0bl15 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b15c710 l0bl15 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b15c711 l0bl15 vdd x711 x711b CELLD r1=10000e3 r0=900e3
xl0b15c712 l0bl15 vdd x712 x712b CELLD r1=10000e3 r0=900e3
xl0b15c713 l0bl15 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b15c714 l0bl15 vdd x714 x714b CELLD r1=10000e3 r0=900e3
xl0b15c715 l0bl15 vdd x715 x715b CELLD r1=10000e3 r0=900e3
xl0b15c716 l0bl15 vdd x716 x716b CELLD r1=10000e3 r0=900e3
xl0b15c717 l0bl15 vdd x717 x717b CELLD r1=10000e3 r0=900e3
xl0b15c718 l0bl15 vdd x718 x718b CELLD r1=10000e3 r0=900e3
xl0b15c719 l0bl15 vdd x719 x719b CELLD r1=900e3 r0=10000e3
xl0b15c720 l0bl15 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b15c721 l0bl15 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b15c722 l0bl15 vdd x722 x722b CELLD r1=10000e3 r0=900e3
xl0b15c723 l0bl15 vdd x723 x723b CELLD r1=900e3 r0=10000e3
xl0b15c724 l0bl15 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b15c725 l0bl15 vdd x725 x725b CELLD r1=900e3 r0=10000e3
xl0b15c726 l0bl15 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b15c727 l0bl15 vdd x727 x727b CELLD r1=10000e3 r0=900e3
xl0b15c728 l0bl15 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b15c729 l0bl15 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b15c730 l0bl15 vdd x730 x730b CELLD r1=900e3 r0=10000e3
xl0b15c731 l0bl15 vdd x731 x731b CELLD r1=900e3 r0=10000e3
xl0b15c732 l0bl15 vdd x732 x732b CELLD r1=10000e3 r0=900e3
xl0b15c733 l0bl15 vdd x733 x733b CELLD r1=10000e3 r0=900e3
xl0b15c734 l0bl15 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b15c735 l0bl15 vdd x735 x735b CELLD r1=10000e3 r0=900e3
xl0b15c736 l0bl15 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b15c737 l0bl15 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b15c738 l0bl15 vdd x738 x738b CELLD r1=10000e3 r0=900e3
xl0b15c739 l0bl15 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b15c740 l0bl15 vdd x740 x740b CELLD r1=10000e3 r0=900e3
xl0b15c741 l0bl15 vdd x741 x741b CELLD r1=10000e3 r0=900e3
xl0b15c742 l0bl15 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b15c743 l0bl15 vdd x743 x743b CELLD r1=10000e3 r0=900e3
xl0b15c744 l0bl15 vdd x744 x744b CELLD r1=10000e3 r0=900e3
xl0b15c745 l0bl15 vdd x745 x745b CELLD r1=10000e3 r0=900e3
xl0b15c746 l0bl15 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b15c747 l0bl15 vdd x747 x747b CELLD r1=900e3 r0=10000e3
xl0b15c748 l0bl15 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b15c749 l0bl15 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b15c750 l0bl15 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b15c751 l0bl15 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b15c752 l0bl15 vdd x752 x752b CELLD r1=900e3 r0=10000e3
xl0b15c753 l0bl15 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b15c754 l0bl15 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b15c755 l0bl15 vdd x755 x755b CELLD r1=900e3 r0=10000e3
xl0b15c756 l0bl15 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b15c757 l0bl15 vdd x757 x757b CELLD r1=10000e3 r0=900e3
xl0b15c758 l0bl15 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b15c759 l0bl15 vdd x759 x759b CELLD r1=900e3 r0=10000e3
xl0b15c760 l0bl15 vdd x760 x760b CELLD r1=900e3 r0=10000e3
xl0b15c761 l0bl15 vdd x761 x761b CELLD r1=900e3 r0=10000e3
xl0b15c762 l0bl15 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b15c763 l0bl15 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b15c764 l0bl15 vdd x764 x764b CELLD r1=10000e3 r0=900e3
xl0b15c765 l0bl15 vdd x765 x765b CELLD r1=10000e3 r0=900e3
xl0b15c766 l0bl15 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b15c767 l0bl15 vdd x767 x767b CELLD r1=10000e3 r0=900e3
xl0b15c768 l0bl15 vdd x768 x768b CELLD r1=10000e3 r0=900e3
xl0b15c769 l0bl15 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b15c770 l0bl15 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b15c771 l0bl15 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b15c772 l0bl15 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b15c773 l0bl15 vdd x773 x773b CELLD r1=10000e3 r0=900e3
xl0b15c774 l0bl15 vdd x774 x774b CELLD r1=10000e3 r0=900e3
xl0b15c775 l0bl15 vdd x775 x775b CELLD r1=10000e3 r0=900e3
xl0b15c776 l0bl15 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b15c777 l0bl15 vdd x777 x777b CELLD r1=900e3 r0=10000e3
xl0b15c778 l0bl15 vdd x778 x778b CELLD r1=900e3 r0=10000e3
xl0b15c779 l0bl15 vdd x779 x779b CELLD r1=900e3 r0=10000e3
xl0b15c780 l0bl15 vdd x780 x780b CELLD r1=900e3 r0=10000e3
xl0b15c781 l0bl15 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b15c782 l0bl15 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b15c783 l0bl15 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b16c0 l0bl16 vdd x0 x0b CELLD r1=10000e3 r0=900e3
xl0b16c1 l0bl16 vdd x1 x1b CELLD r1=10000e3 r0=900e3
xl0b16c2 l0bl16 vdd x2 x2b CELLD r1=10000e3 r0=900e3
xl0b16c3 l0bl16 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b16c4 l0bl16 vdd x4 x4b CELLD r1=900e3 r0=10000e3
xl0b16c5 l0bl16 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b16c6 l0bl16 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b16c7 l0bl16 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b16c8 l0bl16 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b16c9 l0bl16 vdd x9 x9b CELLD r1=10000e3 r0=900e3
xl0b16c10 l0bl16 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b16c11 l0bl16 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b16c12 l0bl16 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b16c13 l0bl16 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b16c14 l0bl16 vdd x14 x14b CELLD r1=10000e3 r0=900e3
xl0b16c15 l0bl16 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b16c16 l0bl16 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b16c17 l0bl16 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b16c18 l0bl16 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b16c19 l0bl16 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b16c20 l0bl16 vdd x20 x20b CELLD r1=900e3 r0=10000e3
xl0b16c21 l0bl16 vdd x21 x21b CELLD r1=10000e3 r0=900e3
xl0b16c22 l0bl16 vdd x22 x22b CELLD r1=10000e3 r0=900e3
xl0b16c23 l0bl16 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b16c24 l0bl16 vdd x24 x24b CELLD r1=900e3 r0=10000e3
xl0b16c25 l0bl16 vdd x25 x25b CELLD r1=10000e3 r0=900e3
xl0b16c26 l0bl16 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b16c27 l0bl16 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b16c28 l0bl16 vdd x28 x28b CELLD r1=10000e3 r0=900e3
xl0b16c29 l0bl16 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b16c30 l0bl16 vdd x30 x30b CELLD r1=900e3 r0=10000e3
xl0b16c31 l0bl16 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b16c32 l0bl16 vdd x32 x32b CELLD r1=10000e3 r0=900e3
xl0b16c33 l0bl16 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b16c34 l0bl16 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b16c35 l0bl16 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b16c36 l0bl16 vdd x36 x36b CELLD r1=10000e3 r0=900e3
xl0b16c37 l0bl16 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b16c38 l0bl16 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b16c39 l0bl16 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b16c40 l0bl16 vdd x40 x40b CELLD r1=900e3 r0=10000e3
xl0b16c41 l0bl16 vdd x41 x41b CELLD r1=10000e3 r0=900e3
xl0b16c42 l0bl16 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b16c43 l0bl16 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b16c44 l0bl16 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b16c45 l0bl16 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b16c46 l0bl16 vdd x46 x46b CELLD r1=10000e3 r0=900e3
xl0b16c47 l0bl16 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b16c48 l0bl16 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b16c49 l0bl16 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b16c50 l0bl16 vdd x50 x50b CELLD r1=10000e3 r0=900e3
xl0b16c51 l0bl16 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b16c52 l0bl16 vdd x52 x52b CELLD r1=10000e3 r0=900e3
xl0b16c53 l0bl16 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b16c54 l0bl16 vdd x54 x54b CELLD r1=10000e3 r0=900e3
xl0b16c55 l0bl16 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b16c56 l0bl16 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b16c57 l0bl16 vdd x57 x57b CELLD r1=10000e3 r0=900e3
xl0b16c58 l0bl16 vdd x58 x58b CELLD r1=900e3 r0=10000e3
xl0b16c59 l0bl16 vdd x59 x59b CELLD r1=10000e3 r0=900e3
xl0b16c60 l0bl16 vdd x60 x60b CELLD r1=10000e3 r0=900e3
xl0b16c61 l0bl16 vdd x61 x61b CELLD r1=10000e3 r0=900e3
xl0b16c62 l0bl16 vdd x62 x62b CELLD r1=10000e3 r0=900e3
xl0b16c63 l0bl16 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b16c64 l0bl16 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b16c65 l0bl16 vdd x65 x65b CELLD r1=10000e3 r0=900e3
xl0b16c66 l0bl16 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b16c67 l0bl16 vdd x67 x67b CELLD r1=10000e3 r0=900e3
xl0b16c68 l0bl16 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b16c69 l0bl16 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b16c70 l0bl16 vdd x70 x70b CELLD r1=10000e3 r0=900e3
xl0b16c71 l0bl16 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b16c72 l0bl16 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b16c73 l0bl16 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b16c74 l0bl16 vdd x74 x74b CELLD r1=10000e3 r0=900e3
xl0b16c75 l0bl16 vdd x75 x75b CELLD r1=10000e3 r0=900e3
xl0b16c76 l0bl16 vdd x76 x76b CELLD r1=10000e3 r0=900e3
xl0b16c77 l0bl16 vdd x77 x77b CELLD r1=10000e3 r0=900e3
xl0b16c78 l0bl16 vdd x78 x78b CELLD r1=10000e3 r0=900e3
xl0b16c79 l0bl16 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b16c80 l0bl16 vdd x80 x80b CELLD r1=10000e3 r0=900e3
xl0b16c81 l0bl16 vdd x81 x81b CELLD r1=10000e3 r0=900e3
xl0b16c82 l0bl16 vdd x82 x82b CELLD r1=10000e3 r0=900e3
xl0b16c83 l0bl16 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b16c84 l0bl16 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b16c85 l0bl16 vdd x85 x85b CELLD r1=10000e3 r0=900e3
xl0b16c86 l0bl16 vdd x86 x86b CELLD r1=900e3 r0=10000e3
xl0b16c87 l0bl16 vdd x87 x87b CELLD r1=10000e3 r0=900e3
xl0b16c88 l0bl16 vdd x88 x88b CELLD r1=10000e3 r0=900e3
xl0b16c89 l0bl16 vdd x89 x89b CELLD r1=900e3 r0=10000e3
xl0b16c90 l0bl16 vdd x90 x90b CELLD r1=10000e3 r0=900e3
xl0b16c91 l0bl16 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b16c92 l0bl16 vdd x92 x92b CELLD r1=900e3 r0=10000e3
xl0b16c93 l0bl16 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b16c94 l0bl16 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b16c95 l0bl16 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b16c96 l0bl16 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b16c97 l0bl16 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b16c98 l0bl16 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b16c99 l0bl16 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b16c100 l0bl16 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b16c101 l0bl16 vdd x101 x101b CELLD r1=900e3 r0=10000e3
xl0b16c102 l0bl16 vdd x102 x102b CELLD r1=10000e3 r0=900e3
xl0b16c103 l0bl16 vdd x103 x103b CELLD r1=10000e3 r0=900e3
xl0b16c104 l0bl16 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b16c105 l0bl16 vdd x105 x105b CELLD r1=10000e3 r0=900e3
xl0b16c106 l0bl16 vdd x106 x106b CELLD r1=10000e3 r0=900e3
xl0b16c107 l0bl16 vdd x107 x107b CELLD r1=10000e3 r0=900e3
xl0b16c108 l0bl16 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b16c109 l0bl16 vdd x109 x109b CELLD r1=10000e3 r0=900e3
xl0b16c110 l0bl16 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b16c111 l0bl16 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b16c112 l0bl16 vdd x112 x112b CELLD r1=10000e3 r0=900e3
xl0b16c113 l0bl16 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b16c114 l0bl16 vdd x114 x114b CELLD r1=10000e3 r0=900e3
xl0b16c115 l0bl16 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b16c116 l0bl16 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b16c117 l0bl16 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b16c118 l0bl16 vdd x118 x118b CELLD r1=10000e3 r0=900e3
xl0b16c119 l0bl16 vdd x119 x119b CELLD r1=10000e3 r0=900e3
xl0b16c120 l0bl16 vdd x120 x120b CELLD r1=900e3 r0=10000e3
xl0b16c121 l0bl16 vdd x121 x121b CELLD r1=900e3 r0=10000e3
xl0b16c122 l0bl16 vdd x122 x122b CELLD r1=900e3 r0=10000e3
xl0b16c123 l0bl16 vdd x123 x123b CELLD r1=900e3 r0=10000e3
xl0b16c124 l0bl16 vdd x124 x124b CELLD r1=900e3 r0=10000e3
xl0b16c125 l0bl16 vdd x125 x125b CELLD r1=900e3 r0=10000e3
xl0b16c126 l0bl16 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b16c127 l0bl16 vdd x127 x127b CELLD r1=900e3 r0=10000e3
xl0b16c128 l0bl16 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b16c129 l0bl16 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b16c130 l0bl16 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b16c131 l0bl16 vdd x131 x131b CELLD r1=10000e3 r0=900e3
xl0b16c132 l0bl16 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b16c133 l0bl16 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b16c134 l0bl16 vdd x134 x134b CELLD r1=10000e3 r0=900e3
xl0b16c135 l0bl16 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b16c136 l0bl16 vdd x136 x136b CELLD r1=900e3 r0=10000e3
xl0b16c137 l0bl16 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b16c138 l0bl16 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b16c139 l0bl16 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b16c140 l0bl16 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b16c141 l0bl16 vdd x141 x141b CELLD r1=10000e3 r0=900e3
xl0b16c142 l0bl16 vdd x142 x142b CELLD r1=900e3 r0=10000e3
xl0b16c143 l0bl16 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b16c144 l0bl16 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b16c145 l0bl16 vdd x145 x145b CELLD r1=900e3 r0=10000e3
xl0b16c146 l0bl16 vdd x146 x146b CELLD r1=900e3 r0=10000e3
xl0b16c147 l0bl16 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b16c148 l0bl16 vdd x148 x148b CELLD r1=900e3 r0=10000e3
xl0b16c149 l0bl16 vdd x149 x149b CELLD r1=900e3 r0=10000e3
xl0b16c150 l0bl16 vdd x150 x150b CELLD r1=900e3 r0=10000e3
xl0b16c151 l0bl16 vdd x151 x151b CELLD r1=900e3 r0=10000e3
xl0b16c152 l0bl16 vdd x152 x152b CELLD r1=900e3 r0=10000e3
xl0b16c153 l0bl16 vdd x153 x153b CELLD r1=900e3 r0=10000e3
xl0b16c154 l0bl16 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b16c155 l0bl16 vdd x155 x155b CELLD r1=900e3 r0=10000e3
xl0b16c156 l0bl16 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b16c157 l0bl16 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b16c158 l0bl16 vdd x158 x158b CELLD r1=10000e3 r0=900e3
xl0b16c159 l0bl16 vdd x159 x159b CELLD r1=10000e3 r0=900e3
xl0b16c160 l0bl16 vdd x160 x160b CELLD r1=10000e3 r0=900e3
xl0b16c161 l0bl16 vdd x161 x161b CELLD r1=10000e3 r0=900e3
xl0b16c162 l0bl16 vdd x162 x162b CELLD r1=10000e3 r0=900e3
xl0b16c163 l0bl16 vdd x163 x163b CELLD r1=10000e3 r0=900e3
xl0b16c164 l0bl16 vdd x164 x164b CELLD r1=10000e3 r0=900e3
xl0b16c165 l0bl16 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b16c166 l0bl16 vdd x166 x166b CELLD r1=10000e3 r0=900e3
xl0b16c167 l0bl16 vdd x167 x167b CELLD r1=10000e3 r0=900e3
xl0b16c168 l0bl16 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b16c169 l0bl16 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b16c170 l0bl16 vdd x170 x170b CELLD r1=10000e3 r0=900e3
xl0b16c171 l0bl16 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b16c172 l0bl16 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b16c173 l0bl16 vdd x173 x173b CELLD r1=10000e3 r0=900e3
xl0b16c174 l0bl16 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b16c175 l0bl16 vdd x175 x175b CELLD r1=900e3 r0=10000e3
xl0b16c176 l0bl16 vdd x176 x176b CELLD r1=900e3 r0=10000e3
xl0b16c177 l0bl16 vdd x177 x177b CELLD r1=900e3 r0=10000e3
xl0b16c178 l0bl16 vdd x178 x178b CELLD r1=900e3 r0=10000e3
xl0b16c179 l0bl16 vdd x179 x179b CELLD r1=900e3 r0=10000e3
xl0b16c180 l0bl16 vdd x180 x180b CELLD r1=900e3 r0=10000e3
xl0b16c181 l0bl16 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b16c182 l0bl16 vdd x182 x182b CELLD r1=900e3 r0=10000e3
xl0b16c183 l0bl16 vdd x183 x183b CELLD r1=900e3 r0=10000e3
xl0b16c184 l0bl16 vdd x184 x184b CELLD r1=900e3 r0=10000e3
xl0b16c185 l0bl16 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b16c186 l0bl16 vdd x186 x186b CELLD r1=10000e3 r0=900e3
xl0b16c187 l0bl16 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b16c188 l0bl16 vdd x188 x188b CELLD r1=10000e3 r0=900e3
xl0b16c189 l0bl16 vdd x189 x189b CELLD r1=10000e3 r0=900e3
xl0b16c190 l0bl16 vdd x190 x190b CELLD r1=10000e3 r0=900e3
xl0b16c191 l0bl16 vdd x191 x191b CELLD r1=10000e3 r0=900e3
xl0b16c192 l0bl16 vdd x192 x192b CELLD r1=10000e3 r0=900e3
xl0b16c193 l0bl16 vdd x193 x193b CELLD r1=900e3 r0=10000e3
xl0b16c194 l0bl16 vdd x194 x194b CELLD r1=10000e3 r0=900e3
xl0b16c195 l0bl16 vdd x195 x195b CELLD r1=10000e3 r0=900e3
xl0b16c196 l0bl16 vdd x196 x196b CELLD r1=10000e3 r0=900e3
xl0b16c197 l0bl16 vdd x197 x197b CELLD r1=10000e3 r0=900e3
xl0b16c198 l0bl16 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b16c199 l0bl16 vdd x199 x199b CELLD r1=10000e3 r0=900e3
xl0b16c200 l0bl16 vdd x200 x200b CELLD r1=10000e3 r0=900e3
xl0b16c201 l0bl16 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b16c202 l0bl16 vdd x202 x202b CELLD r1=900e3 r0=10000e3
xl0b16c203 l0bl16 vdd x203 x203b CELLD r1=900e3 r0=10000e3
xl0b16c204 l0bl16 vdd x204 x204b CELLD r1=900e3 r0=10000e3
xl0b16c205 l0bl16 vdd x205 x205b CELLD r1=900e3 r0=10000e3
xl0b16c206 l0bl16 vdd x206 x206b CELLD r1=900e3 r0=10000e3
xl0b16c207 l0bl16 vdd x207 x207b CELLD r1=900e3 r0=10000e3
xl0b16c208 l0bl16 vdd x208 x208b CELLD r1=900e3 r0=10000e3
xl0b16c209 l0bl16 vdd x209 x209b CELLD r1=900e3 r0=10000e3
xl0b16c210 l0bl16 vdd x210 x210b CELLD r1=900e3 r0=10000e3
xl0b16c211 l0bl16 vdd x211 x211b CELLD r1=900e3 r0=10000e3
xl0b16c212 l0bl16 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b16c213 l0bl16 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b16c214 l0bl16 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b16c215 l0bl16 vdd x215 x215b CELLD r1=900e3 r0=10000e3
xl0b16c216 l0bl16 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b16c217 l0bl16 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b16c218 l0bl16 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b16c219 l0bl16 vdd x219 x219b CELLD r1=10000e3 r0=900e3
xl0b16c220 l0bl16 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b16c221 l0bl16 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b16c222 l0bl16 vdd x222 x222b CELLD r1=10000e3 r0=900e3
xl0b16c223 l0bl16 vdd x223 x223b CELLD r1=900e3 r0=10000e3
xl0b16c224 l0bl16 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b16c225 l0bl16 vdd x225 x225b CELLD r1=900e3 r0=10000e3
xl0b16c226 l0bl16 vdd x226 x226b CELLD r1=900e3 r0=10000e3
xl0b16c227 l0bl16 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b16c228 l0bl16 vdd x228 x228b CELLD r1=900e3 r0=10000e3
xl0b16c229 l0bl16 vdd x229 x229b CELLD r1=10000e3 r0=900e3
xl0b16c230 l0bl16 vdd x230 x230b CELLD r1=900e3 r0=10000e3
xl0b16c231 l0bl16 vdd x231 x231b CELLD r1=900e3 r0=10000e3
xl0b16c232 l0bl16 vdd x232 x232b CELLD r1=900e3 r0=10000e3
xl0b16c233 l0bl16 vdd x233 x233b CELLD r1=900e3 r0=10000e3
xl0b16c234 l0bl16 vdd x234 x234b CELLD r1=900e3 r0=10000e3
xl0b16c235 l0bl16 vdd x235 x235b CELLD r1=900e3 r0=10000e3
xl0b16c236 l0bl16 vdd x236 x236b CELLD r1=900e3 r0=10000e3
xl0b16c237 l0bl16 vdd x237 x237b CELLD r1=900e3 r0=10000e3
xl0b16c238 l0bl16 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b16c239 l0bl16 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b16c240 l0bl16 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b16c241 l0bl16 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b16c242 l0bl16 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b16c243 l0bl16 vdd x243 x243b CELLD r1=900e3 r0=10000e3
xl0b16c244 l0bl16 vdd x244 x244b CELLD r1=900e3 r0=10000e3
xl0b16c245 l0bl16 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b16c246 l0bl16 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b16c247 l0bl16 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b16c248 l0bl16 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b16c249 l0bl16 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b16c250 l0bl16 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b16c251 l0bl16 vdd x251 x251b CELLD r1=900e3 r0=10000e3
xl0b16c252 l0bl16 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b16c253 l0bl16 vdd x253 x253b CELLD r1=10000e3 r0=900e3
xl0b16c254 l0bl16 vdd x254 x254b CELLD r1=900e3 r0=10000e3
xl0b16c255 l0bl16 vdd x255 x255b CELLD r1=900e3 r0=10000e3
xl0b16c256 l0bl16 vdd x256 x256b CELLD r1=10000e3 r0=900e3
xl0b16c257 l0bl16 vdd x257 x257b CELLD r1=900e3 r0=10000e3
xl0b16c258 l0bl16 vdd x258 x258b CELLD r1=900e3 r0=10000e3
xl0b16c259 l0bl16 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b16c260 l0bl16 vdd x260 x260b CELLD r1=900e3 r0=10000e3
xl0b16c261 l0bl16 vdd x261 x261b CELLD r1=900e3 r0=10000e3
xl0b16c262 l0bl16 vdd x262 x262b CELLD r1=900e3 r0=10000e3
xl0b16c263 l0bl16 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b16c264 l0bl16 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b16c265 l0bl16 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b16c266 l0bl16 vdd x266 x266b CELLD r1=900e3 r0=10000e3
xl0b16c267 l0bl16 vdd x267 x267b CELLD r1=900e3 r0=10000e3
xl0b16c268 l0bl16 vdd x268 x268b CELLD r1=900e3 r0=10000e3
xl0b16c269 l0bl16 vdd x269 x269b CELLD r1=900e3 r0=10000e3
xl0b16c270 l0bl16 vdd x270 x270b CELLD r1=900e3 r0=10000e3
xl0b16c271 l0bl16 vdd x271 x271b CELLD r1=900e3 r0=10000e3
xl0b16c272 l0bl16 vdd x272 x272b CELLD r1=900e3 r0=10000e3
xl0b16c273 l0bl16 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b16c274 l0bl16 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b16c275 l0bl16 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b16c276 l0bl16 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b16c277 l0bl16 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b16c278 l0bl16 vdd x278 x278b CELLD r1=900e3 r0=10000e3
xl0b16c279 l0bl16 vdd x279 x279b CELLD r1=10000e3 r0=900e3
xl0b16c280 l0bl16 vdd x280 x280b CELLD r1=10000e3 r0=900e3
xl0b16c281 l0bl16 vdd x281 x281b CELLD r1=900e3 r0=10000e3
xl0b16c282 l0bl16 vdd x282 x282b CELLD r1=900e3 r0=10000e3
xl0b16c283 l0bl16 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b16c284 l0bl16 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b16c285 l0bl16 vdd x285 x285b CELLD r1=900e3 r0=10000e3
xl0b16c286 l0bl16 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b16c287 l0bl16 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b16c288 l0bl16 vdd x288 x288b CELLD r1=900e3 r0=10000e3
xl0b16c289 l0bl16 vdd x289 x289b CELLD r1=900e3 r0=10000e3
xl0b16c290 l0bl16 vdd x290 x290b CELLD r1=10000e3 r0=900e3
xl0b16c291 l0bl16 vdd x291 x291b CELLD r1=10000e3 r0=900e3
xl0b16c292 l0bl16 vdd x292 x292b CELLD r1=10000e3 r0=900e3
xl0b16c293 l0bl16 vdd x293 x293b CELLD r1=10000e3 r0=900e3
xl0b16c294 l0bl16 vdd x294 x294b CELLD r1=10000e3 r0=900e3
xl0b16c295 l0bl16 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b16c296 l0bl16 vdd x296 x296b CELLD r1=900e3 r0=10000e3
xl0b16c297 l0bl16 vdd x297 x297b CELLD r1=900e3 r0=10000e3
xl0b16c298 l0bl16 vdd x298 x298b CELLD r1=900e3 r0=10000e3
xl0b16c299 l0bl16 vdd x299 x299b CELLD r1=900e3 r0=10000e3
xl0b16c300 l0bl16 vdd x300 x300b CELLD r1=900e3 r0=10000e3
xl0b16c301 l0bl16 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b16c302 l0bl16 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b16c303 l0bl16 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b16c304 l0bl16 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b16c305 l0bl16 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b16c306 l0bl16 vdd x306 x306b CELLD r1=10000e3 r0=900e3
xl0b16c307 l0bl16 vdd x307 x307b CELLD r1=900e3 r0=10000e3
xl0b16c308 l0bl16 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b16c309 l0bl16 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b16c310 l0bl16 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b16c311 l0bl16 vdd x311 x311b CELLD r1=900e3 r0=10000e3
xl0b16c312 l0bl16 vdd x312 x312b CELLD r1=900e3 r0=10000e3
xl0b16c313 l0bl16 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b16c314 l0bl16 vdd x314 x314b CELLD r1=900e3 r0=10000e3
xl0b16c315 l0bl16 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b16c316 l0bl16 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b16c317 l0bl16 vdd x317 x317b CELLD r1=10000e3 r0=900e3
xl0b16c318 l0bl16 vdd x318 x318b CELLD r1=10000e3 r0=900e3
xl0b16c319 l0bl16 vdd x319 x319b CELLD r1=10000e3 r0=900e3
xl0b16c320 l0bl16 vdd x320 x320b CELLD r1=10000e3 r0=900e3
xl0b16c321 l0bl16 vdd x321 x321b CELLD r1=10000e3 r0=900e3
xl0b16c322 l0bl16 vdd x322 x322b CELLD r1=10000e3 r0=900e3
xl0b16c323 l0bl16 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b16c324 l0bl16 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b16c325 l0bl16 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b16c326 l0bl16 vdd x326 x326b CELLD r1=900e3 r0=10000e3
xl0b16c327 l0bl16 vdd x327 x327b CELLD r1=900e3 r0=10000e3
xl0b16c328 l0bl16 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b16c329 l0bl16 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b16c330 l0bl16 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b16c331 l0bl16 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b16c332 l0bl16 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b16c333 l0bl16 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b16c334 l0bl16 vdd x334 x334b CELLD r1=10000e3 r0=900e3
xl0b16c335 l0bl16 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b16c336 l0bl16 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b16c337 l0bl16 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b16c338 l0bl16 vdd x338 x338b CELLD r1=900e3 r0=10000e3
xl0b16c339 l0bl16 vdd x339 x339b CELLD r1=900e3 r0=10000e3
xl0b16c340 l0bl16 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b16c341 l0bl16 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b16c342 l0bl16 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b16c343 l0bl16 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b16c344 l0bl16 vdd x344 x344b CELLD r1=10000e3 r0=900e3
xl0b16c345 l0bl16 vdd x345 x345b CELLD r1=10000e3 r0=900e3
xl0b16c346 l0bl16 vdd x346 x346b CELLD r1=10000e3 r0=900e3
xl0b16c347 l0bl16 vdd x347 x347b CELLD r1=10000e3 r0=900e3
xl0b16c348 l0bl16 vdd x348 x348b CELLD r1=10000e3 r0=900e3
xl0b16c349 l0bl16 vdd x349 x349b CELLD r1=10000e3 r0=900e3
xl0b16c350 l0bl16 vdd x350 x350b CELLD r1=10000e3 r0=900e3
xl0b16c351 l0bl16 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b16c352 l0bl16 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b16c353 l0bl16 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b16c354 l0bl16 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b16c355 l0bl16 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b16c356 l0bl16 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b16c357 l0bl16 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b16c358 l0bl16 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b16c359 l0bl16 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b16c360 l0bl16 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b16c361 l0bl16 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b16c362 l0bl16 vdd x362 x362b CELLD r1=10000e3 r0=900e3
xl0b16c363 l0bl16 vdd x363 x363b CELLD r1=10000e3 r0=900e3
xl0b16c364 l0bl16 vdd x364 x364b CELLD r1=900e3 r0=10000e3
xl0b16c365 l0bl16 vdd x365 x365b CELLD r1=10000e3 r0=900e3
xl0b16c366 l0bl16 vdd x366 x366b CELLD r1=10000e3 r0=900e3
xl0b16c367 l0bl16 vdd x367 x367b CELLD r1=900e3 r0=10000e3
xl0b16c368 l0bl16 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b16c369 l0bl16 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b16c370 l0bl16 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b16c371 l0bl16 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b16c372 l0bl16 vdd x372 x372b CELLD r1=10000e3 r0=900e3
xl0b16c373 l0bl16 vdd x373 x373b CELLD r1=10000e3 r0=900e3
xl0b16c374 l0bl16 vdd x374 x374b CELLD r1=10000e3 r0=900e3
xl0b16c375 l0bl16 vdd x375 x375b CELLD r1=10000e3 r0=900e3
xl0b16c376 l0bl16 vdd x376 x376b CELLD r1=10000e3 r0=900e3
xl0b16c377 l0bl16 vdd x377 x377b CELLD r1=10000e3 r0=900e3
xl0b16c378 l0bl16 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b16c379 l0bl16 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b16c380 l0bl16 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b16c381 l0bl16 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b16c382 l0bl16 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b16c383 l0bl16 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b16c384 l0bl16 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b16c385 l0bl16 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b16c386 l0bl16 vdd x386 x386b CELLD r1=10000e3 r0=900e3
xl0b16c387 l0bl16 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b16c388 l0bl16 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b16c389 l0bl16 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b16c390 l0bl16 vdd x390 x390b CELLD r1=900e3 r0=10000e3
xl0b16c391 l0bl16 vdd x391 x391b CELLD r1=900e3 r0=10000e3
xl0b16c392 l0bl16 vdd x392 x392b CELLD r1=10000e3 r0=900e3
xl0b16c393 l0bl16 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b16c394 l0bl16 vdd x394 x394b CELLD r1=10000e3 r0=900e3
xl0b16c395 l0bl16 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b16c396 l0bl16 vdd x396 x396b CELLD r1=900e3 r0=10000e3
xl0b16c397 l0bl16 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b16c398 l0bl16 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b16c399 l0bl16 vdd x399 x399b CELLD r1=10000e3 r0=900e3
xl0b16c400 l0bl16 vdd x400 x400b CELLD r1=10000e3 r0=900e3
xl0b16c401 l0bl16 vdd x401 x401b CELLD r1=10000e3 r0=900e3
xl0b16c402 l0bl16 vdd x402 x402b CELLD r1=10000e3 r0=900e3
xl0b16c403 l0bl16 vdd x403 x403b CELLD r1=10000e3 r0=900e3
xl0b16c404 l0bl16 vdd x404 x404b CELLD r1=10000e3 r0=900e3
xl0b16c405 l0bl16 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b16c406 l0bl16 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b16c407 l0bl16 vdd x407 x407b CELLD r1=900e3 r0=10000e3
xl0b16c408 l0bl16 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b16c409 l0bl16 vdd x409 x409b CELLD r1=10000e3 r0=900e3
xl0b16c410 l0bl16 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b16c411 l0bl16 vdd x411 x411b CELLD r1=10000e3 r0=900e3
xl0b16c412 l0bl16 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b16c413 l0bl16 vdd x413 x413b CELLD r1=10000e3 r0=900e3
xl0b16c414 l0bl16 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b16c415 l0bl16 vdd x415 x415b CELLD r1=10000e3 r0=900e3
xl0b16c416 l0bl16 vdd x416 x416b CELLD r1=900e3 r0=10000e3
xl0b16c417 l0bl16 vdd x417 x417b CELLD r1=900e3 r0=10000e3
xl0b16c418 l0bl16 vdd x418 x418b CELLD r1=900e3 r0=10000e3
xl0b16c419 l0bl16 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b16c420 l0bl16 vdd x420 x420b CELLD r1=900e3 r0=10000e3
xl0b16c421 l0bl16 vdd x421 x421b CELLD r1=900e3 r0=10000e3
xl0b16c422 l0bl16 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b16c423 l0bl16 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b16c424 l0bl16 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b16c425 l0bl16 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b16c426 l0bl16 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b16c427 l0bl16 vdd x427 x427b CELLD r1=10000e3 r0=900e3
xl0b16c428 l0bl16 vdd x428 x428b CELLD r1=10000e3 r0=900e3
xl0b16c429 l0bl16 vdd x429 x429b CELLD r1=10000e3 r0=900e3
xl0b16c430 l0bl16 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b16c431 l0bl16 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b16c432 l0bl16 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b16c433 l0bl16 vdd x433 x433b CELLD r1=900e3 r0=10000e3
xl0b16c434 l0bl16 vdd x434 x434b CELLD r1=900e3 r0=10000e3
xl0b16c435 l0bl16 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b16c436 l0bl16 vdd x436 x436b CELLD r1=10000e3 r0=900e3
xl0b16c437 l0bl16 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b16c438 l0bl16 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b16c439 l0bl16 vdd x439 x439b CELLD r1=10000e3 r0=900e3
xl0b16c440 l0bl16 vdd x440 x440b CELLD r1=10000e3 r0=900e3
xl0b16c441 l0bl16 vdd x441 x441b CELLD r1=10000e3 r0=900e3
xl0b16c442 l0bl16 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b16c443 l0bl16 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b16c444 l0bl16 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b16c445 l0bl16 vdd x445 x445b CELLD r1=900e3 r0=10000e3
xl0b16c446 l0bl16 vdd x446 x446b CELLD r1=900e3 r0=10000e3
xl0b16c447 l0bl16 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b16c448 l0bl16 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b16c449 l0bl16 vdd x449 x449b CELLD r1=10000e3 r0=900e3
xl0b16c450 l0bl16 vdd x450 x450b CELLD r1=10000e3 r0=900e3
xl0b16c451 l0bl16 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b16c452 l0bl16 vdd x452 x452b CELLD r1=900e3 r0=10000e3
xl0b16c453 l0bl16 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b16c454 l0bl16 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b16c455 l0bl16 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b16c456 l0bl16 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b16c457 l0bl16 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b16c458 l0bl16 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b16c459 l0bl16 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b16c460 l0bl16 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b16c461 l0bl16 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b16c462 l0bl16 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b16c463 l0bl16 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b16c464 l0bl16 vdd x464 x464b CELLD r1=10000e3 r0=900e3
xl0b16c465 l0bl16 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b16c466 l0bl16 vdd x466 x466b CELLD r1=10000e3 r0=900e3
xl0b16c467 l0bl16 vdd x467 x467b CELLD r1=10000e3 r0=900e3
xl0b16c468 l0bl16 vdd x468 x468b CELLD r1=10000e3 r0=900e3
xl0b16c469 l0bl16 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b16c470 l0bl16 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b16c471 l0bl16 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b16c472 l0bl16 vdd x472 x472b CELLD r1=900e3 r0=10000e3
xl0b16c473 l0bl16 vdd x473 x473b CELLD r1=900e3 r0=10000e3
xl0b16c474 l0bl16 vdd x474 x474b CELLD r1=10000e3 r0=900e3
xl0b16c475 l0bl16 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b16c476 l0bl16 vdd x476 x476b CELLD r1=10000e3 r0=900e3
xl0b16c477 l0bl16 vdd x477 x477b CELLD r1=10000e3 r0=900e3
xl0b16c478 l0bl16 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b16c479 l0bl16 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b16c480 l0bl16 vdd x480 x480b CELLD r1=900e3 r0=10000e3
xl0b16c481 l0bl16 vdd x481 x481b CELLD r1=900e3 r0=10000e3
xl0b16c482 l0bl16 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b16c483 l0bl16 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b16c484 l0bl16 vdd x484 x484b CELLD r1=900e3 r0=10000e3
xl0b16c485 l0bl16 vdd x485 x485b CELLD r1=900e3 r0=10000e3
xl0b16c486 l0bl16 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b16c487 l0bl16 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b16c488 l0bl16 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b16c489 l0bl16 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b16c490 l0bl16 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b16c491 l0bl16 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b16c492 l0bl16 vdd x492 x492b CELLD r1=10000e3 r0=900e3
xl0b16c493 l0bl16 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b16c494 l0bl16 vdd x494 x494b CELLD r1=10000e3 r0=900e3
xl0b16c495 l0bl16 vdd x495 x495b CELLD r1=900e3 r0=10000e3
xl0b16c496 l0bl16 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b16c497 l0bl16 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b16c498 l0bl16 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b16c499 l0bl16 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b16c500 l0bl16 vdd x500 x500b CELLD r1=900e3 r0=10000e3
xl0b16c501 l0bl16 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b16c502 l0bl16 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b16c503 l0bl16 vdd x503 x503b CELLD r1=10000e3 r0=900e3
xl0b16c504 l0bl16 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b16c505 l0bl16 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b16c506 l0bl16 vdd x506 x506b CELLD r1=900e3 r0=10000e3
xl0b16c507 l0bl16 vdd x507 x507b CELLD r1=900e3 r0=10000e3
xl0b16c508 l0bl16 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b16c509 l0bl16 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b16c510 l0bl16 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b16c511 l0bl16 vdd x511 x511b CELLD r1=900e3 r0=10000e3
xl0b16c512 l0bl16 vdd x512 x512b CELLD r1=900e3 r0=10000e3
xl0b16c513 l0bl16 vdd x513 x513b CELLD r1=900e3 r0=10000e3
xl0b16c514 l0bl16 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b16c515 l0bl16 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b16c516 l0bl16 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b16c517 l0bl16 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b16c518 l0bl16 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b16c519 l0bl16 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b16c520 l0bl16 vdd x520 x520b CELLD r1=10000e3 r0=900e3
xl0b16c521 l0bl16 vdd x521 x521b CELLD r1=10000e3 r0=900e3
xl0b16c522 l0bl16 vdd x522 x522b CELLD r1=10000e3 r0=900e3
xl0b16c523 l0bl16 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b16c524 l0bl16 vdd x524 x524b CELLD r1=900e3 r0=10000e3
xl0b16c525 l0bl16 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b16c526 l0bl16 vdd x526 x526b CELLD r1=900e3 r0=10000e3
xl0b16c527 l0bl16 vdd x527 x527b CELLD r1=900e3 r0=10000e3
xl0b16c528 l0bl16 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b16c529 l0bl16 vdd x529 x529b CELLD r1=900e3 r0=10000e3
xl0b16c530 l0bl16 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b16c531 l0bl16 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b16c532 l0bl16 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b16c533 l0bl16 vdd x533 x533b CELLD r1=10000e3 r0=900e3
xl0b16c534 l0bl16 vdd x534 x534b CELLD r1=10000e3 r0=900e3
xl0b16c535 l0bl16 vdd x535 x535b CELLD r1=10000e3 r0=900e3
xl0b16c536 l0bl16 vdd x536 x536b CELLD r1=900e3 r0=10000e3
xl0b16c537 l0bl16 vdd x537 x537b CELLD r1=900e3 r0=10000e3
xl0b16c538 l0bl16 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b16c539 l0bl16 vdd x539 x539b CELLD r1=900e3 r0=10000e3
xl0b16c540 l0bl16 vdd x540 x540b CELLD r1=900e3 r0=10000e3
xl0b16c541 l0bl16 vdd x541 x541b CELLD r1=900e3 r0=10000e3
xl0b16c542 l0bl16 vdd x542 x542b CELLD r1=900e3 r0=10000e3
xl0b16c543 l0bl16 vdd x543 x543b CELLD r1=900e3 r0=10000e3
xl0b16c544 l0bl16 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b16c545 l0bl16 vdd x545 x545b CELLD r1=900e3 r0=10000e3
xl0b16c546 l0bl16 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b16c547 l0bl16 vdd x547 x547b CELLD r1=10000e3 r0=900e3
xl0b16c548 l0bl16 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b16c549 l0bl16 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b16c550 l0bl16 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b16c551 l0bl16 vdd x551 x551b CELLD r1=900e3 r0=10000e3
xl0b16c552 l0bl16 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b16c553 l0bl16 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b16c554 l0bl16 vdd x554 x554b CELLD r1=900e3 r0=10000e3
xl0b16c555 l0bl16 vdd x555 x555b CELLD r1=900e3 r0=10000e3
xl0b16c556 l0bl16 vdd x556 x556b CELLD r1=900e3 r0=10000e3
xl0b16c557 l0bl16 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b16c558 l0bl16 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b16c559 l0bl16 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b16c560 l0bl16 vdd x560 x560b CELLD r1=10000e3 r0=900e3
xl0b16c561 l0bl16 vdd x561 x561b CELLD r1=10000e3 r0=900e3
xl0b16c562 l0bl16 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b16c563 l0bl16 vdd x563 x563b CELLD r1=900e3 r0=10000e3
xl0b16c564 l0bl16 vdd x564 x564b CELLD r1=900e3 r0=10000e3
xl0b16c565 l0bl16 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b16c566 l0bl16 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b16c567 l0bl16 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b16c568 l0bl16 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b16c569 l0bl16 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b16c570 l0bl16 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b16c571 l0bl16 vdd x571 x571b CELLD r1=10000e3 r0=900e3
xl0b16c572 l0bl16 vdd x572 x572b CELLD r1=10000e3 r0=900e3
xl0b16c573 l0bl16 vdd x573 x573b CELLD r1=10000e3 r0=900e3
xl0b16c574 l0bl16 vdd x574 x574b CELLD r1=10000e3 r0=900e3
xl0b16c575 l0bl16 vdd x575 x575b CELLD r1=10000e3 r0=900e3
xl0b16c576 l0bl16 vdd x576 x576b CELLD r1=10000e3 r0=900e3
xl0b16c577 l0bl16 vdd x577 x577b CELLD r1=900e3 r0=10000e3
xl0b16c578 l0bl16 vdd x578 x578b CELLD r1=10000e3 r0=900e3
xl0b16c579 l0bl16 vdd x579 x579b CELLD r1=10000e3 r0=900e3
xl0b16c580 l0bl16 vdd x580 x580b CELLD r1=10000e3 r0=900e3
xl0b16c581 l0bl16 vdd x581 x581b CELLD r1=900e3 r0=10000e3
xl0b16c582 l0bl16 vdd x582 x582b CELLD r1=900e3 r0=10000e3
xl0b16c583 l0bl16 vdd x583 x583b CELLD r1=900e3 r0=10000e3
xl0b16c584 l0bl16 vdd x584 x584b CELLD r1=900e3 r0=10000e3
xl0b16c585 l0bl16 vdd x585 x585b CELLD r1=900e3 r0=10000e3
xl0b16c586 l0bl16 vdd x586 x586b CELLD r1=900e3 r0=10000e3
xl0b16c587 l0bl16 vdd x587 x587b CELLD r1=900e3 r0=10000e3
xl0b16c588 l0bl16 vdd x588 x588b CELLD r1=900e3 r0=10000e3
xl0b16c589 l0bl16 vdd x589 x589b CELLD r1=900e3 r0=10000e3
xl0b16c590 l0bl16 vdd x590 x590b CELLD r1=900e3 r0=10000e3
xl0b16c591 l0bl16 vdd x591 x591b CELLD r1=10000e3 r0=900e3
xl0b16c592 l0bl16 vdd x592 x592b CELLD r1=10000e3 r0=900e3
xl0b16c593 l0bl16 vdd x593 x593b CELLD r1=10000e3 r0=900e3
xl0b16c594 l0bl16 vdd x594 x594b CELLD r1=10000e3 r0=900e3
xl0b16c595 l0bl16 vdd x595 x595b CELLD r1=10000e3 r0=900e3
xl0b16c596 l0bl16 vdd x596 x596b CELLD r1=10000e3 r0=900e3
xl0b16c597 l0bl16 vdd x597 x597b CELLD r1=10000e3 r0=900e3
xl0b16c598 l0bl16 vdd x598 x598b CELLD r1=10000e3 r0=900e3
xl0b16c599 l0bl16 vdd x599 x599b CELLD r1=10000e3 r0=900e3
xl0b16c600 l0bl16 vdd x600 x600b CELLD r1=10000e3 r0=900e3
xl0b16c601 l0bl16 vdd x601 x601b CELLD r1=10000e3 r0=900e3
xl0b16c602 l0bl16 vdd x602 x602b CELLD r1=10000e3 r0=900e3
xl0b16c603 l0bl16 vdd x603 x603b CELLD r1=10000e3 r0=900e3
xl0b16c604 l0bl16 vdd x604 x604b CELLD r1=10000e3 r0=900e3
xl0b16c605 l0bl16 vdd x605 x605b CELLD r1=10000e3 r0=900e3
xl0b16c606 l0bl16 vdd x606 x606b CELLD r1=10000e3 r0=900e3
xl0b16c607 l0bl16 vdd x607 x607b CELLD r1=900e3 r0=10000e3
xl0b16c608 l0bl16 vdd x608 x608b CELLD r1=900e3 r0=10000e3
xl0b16c609 l0bl16 vdd x609 x609b CELLD r1=900e3 r0=10000e3
xl0b16c610 l0bl16 vdd x610 x610b CELLD r1=900e3 r0=10000e3
xl0b16c611 l0bl16 vdd x611 x611b CELLD r1=900e3 r0=10000e3
xl0b16c612 l0bl16 vdd x612 x612b CELLD r1=10000e3 r0=900e3
xl0b16c613 l0bl16 vdd x613 x613b CELLD r1=10000e3 r0=900e3
xl0b16c614 l0bl16 vdd x614 x614b CELLD r1=900e3 r0=10000e3
xl0b16c615 l0bl16 vdd x615 x615b CELLD r1=10000e3 r0=900e3
xl0b16c616 l0bl16 vdd x616 x616b CELLD r1=900e3 r0=10000e3
xl0b16c617 l0bl16 vdd x617 x617b CELLD r1=900e3 r0=10000e3
xl0b16c618 l0bl16 vdd x618 x618b CELLD r1=900e3 r0=10000e3
xl0b16c619 l0bl16 vdd x619 x619b CELLD r1=10000e3 r0=900e3
xl0b16c620 l0bl16 vdd x620 x620b CELLD r1=10000e3 r0=900e3
xl0b16c621 l0bl16 vdd x621 x621b CELLD r1=10000e3 r0=900e3
xl0b16c622 l0bl16 vdd x622 x622b CELLD r1=900e3 r0=10000e3
xl0b16c623 l0bl16 vdd x623 x623b CELLD r1=10000e3 r0=900e3
xl0b16c624 l0bl16 vdd x624 x624b CELLD r1=900e3 r0=10000e3
xl0b16c625 l0bl16 vdd x625 x625b CELLD r1=10000e3 r0=900e3
xl0b16c626 l0bl16 vdd x626 x626b CELLD r1=10000e3 r0=900e3
xl0b16c627 l0bl16 vdd x627 x627b CELLD r1=10000e3 r0=900e3
xl0b16c628 l0bl16 vdd x628 x628b CELLD r1=10000e3 r0=900e3
xl0b16c629 l0bl16 vdd x629 x629b CELLD r1=10000e3 r0=900e3
xl0b16c630 l0bl16 vdd x630 x630b CELLD r1=10000e3 r0=900e3
xl0b16c631 l0bl16 vdd x631 x631b CELLD r1=10000e3 r0=900e3
xl0b16c632 l0bl16 vdd x632 x632b CELLD r1=10000e3 r0=900e3
xl0b16c633 l0bl16 vdd x633 x633b CELLD r1=900e3 r0=10000e3
xl0b16c634 l0bl16 vdd x634 x634b CELLD r1=900e3 r0=10000e3
xl0b16c635 l0bl16 vdd x635 x635b CELLD r1=900e3 r0=10000e3
xl0b16c636 l0bl16 vdd x636 x636b CELLD r1=900e3 r0=10000e3
xl0b16c637 l0bl16 vdd x637 x637b CELLD r1=900e3 r0=10000e3
xl0b16c638 l0bl16 vdd x638 x638b CELLD r1=900e3 r0=10000e3
xl0b16c639 l0bl16 vdd x639 x639b CELLD r1=900e3 r0=10000e3
xl0b16c640 l0bl16 vdd x640 x640b CELLD r1=900e3 r0=10000e3
xl0b16c641 l0bl16 vdd x641 x641b CELLD r1=900e3 r0=10000e3
xl0b16c642 l0bl16 vdd x642 x642b CELLD r1=900e3 r0=10000e3
xl0b16c643 l0bl16 vdd x643 x643b CELLD r1=900e3 r0=10000e3
xl0b16c644 l0bl16 vdd x644 x644b CELLD r1=10000e3 r0=900e3
xl0b16c645 l0bl16 vdd x645 x645b CELLD r1=900e3 r0=10000e3
xl0b16c646 l0bl16 vdd x646 x646b CELLD r1=10000e3 r0=900e3
xl0b16c647 l0bl16 vdd x647 x647b CELLD r1=10000e3 r0=900e3
xl0b16c648 l0bl16 vdd x648 x648b CELLD r1=900e3 r0=10000e3
xl0b16c649 l0bl16 vdd x649 x649b CELLD r1=10000e3 r0=900e3
xl0b16c650 l0bl16 vdd x650 x650b CELLD r1=10000e3 r0=900e3
xl0b16c651 l0bl16 vdd x651 x651b CELLD r1=900e3 r0=10000e3
xl0b16c652 l0bl16 vdd x652 x652b CELLD r1=10000e3 r0=900e3
xl0b16c653 l0bl16 vdd x653 x653b CELLD r1=900e3 r0=10000e3
xl0b16c654 l0bl16 vdd x654 x654b CELLD r1=10000e3 r0=900e3
xl0b16c655 l0bl16 vdd x655 x655b CELLD r1=10000e3 r0=900e3
xl0b16c656 l0bl16 vdd x656 x656b CELLD r1=10000e3 r0=900e3
xl0b16c657 l0bl16 vdd x657 x657b CELLD r1=10000e3 r0=900e3
xl0b16c658 l0bl16 vdd x658 x658b CELLD r1=10000e3 r0=900e3
xl0b16c659 l0bl16 vdd x659 x659b CELLD r1=10000e3 r0=900e3
xl0b16c660 l0bl16 vdd x660 x660b CELLD r1=10000e3 r0=900e3
xl0b16c661 l0bl16 vdd x661 x661b CELLD r1=900e3 r0=10000e3
xl0b16c662 l0bl16 vdd x662 x662b CELLD r1=900e3 r0=10000e3
xl0b16c663 l0bl16 vdd x663 x663b CELLD r1=900e3 r0=10000e3
xl0b16c664 l0bl16 vdd x664 x664b CELLD r1=900e3 r0=10000e3
xl0b16c665 l0bl16 vdd x665 x665b CELLD r1=900e3 r0=10000e3
xl0b16c666 l0bl16 vdd x666 x666b CELLD r1=10000e3 r0=900e3
xl0b16c667 l0bl16 vdd x667 x667b CELLD r1=10000e3 r0=900e3
xl0b16c668 l0bl16 vdd x668 x668b CELLD r1=900e3 r0=10000e3
xl0b16c669 l0bl16 vdd x669 x669b CELLD r1=900e3 r0=10000e3
xl0b16c670 l0bl16 vdd x670 x670b CELLD r1=900e3 r0=10000e3
xl0b16c671 l0bl16 vdd x671 x671b CELLD r1=900e3 r0=10000e3
xl0b16c672 l0bl16 vdd x672 x672b CELLD r1=10000e3 r0=900e3
xl0b16c673 l0bl16 vdd x673 x673b CELLD r1=900e3 r0=10000e3
xl0b16c674 l0bl16 vdd x674 x674b CELLD r1=10000e3 r0=900e3
xl0b16c675 l0bl16 vdd x675 x675b CELLD r1=10000e3 r0=900e3
xl0b16c676 l0bl16 vdd x676 x676b CELLD r1=10000e3 r0=900e3
xl0b16c677 l0bl16 vdd x677 x677b CELLD r1=900e3 r0=10000e3
xl0b16c678 l0bl16 vdd x678 x678b CELLD r1=900e3 r0=10000e3
xl0b16c679 l0bl16 vdd x679 x679b CELLD r1=900e3 r0=10000e3
xl0b16c680 l0bl16 vdd x680 x680b CELLD r1=900e3 r0=10000e3
xl0b16c681 l0bl16 vdd x681 x681b CELLD r1=900e3 r0=10000e3
xl0b16c682 l0bl16 vdd x682 x682b CELLD r1=900e3 r0=10000e3
xl0b16c683 l0bl16 vdd x683 x683b CELLD r1=10000e3 r0=900e3
xl0b16c684 l0bl16 vdd x684 x684b CELLD r1=10000e3 r0=900e3
xl0b16c685 l0bl16 vdd x685 x685b CELLD r1=10000e3 r0=900e3
xl0b16c686 l0bl16 vdd x686 x686b CELLD r1=900e3 r0=10000e3
xl0b16c687 l0bl16 vdd x687 x687b CELLD r1=900e3 r0=10000e3
xl0b16c688 l0bl16 vdd x688 x688b CELLD r1=900e3 r0=10000e3
xl0b16c689 l0bl16 vdd x689 x689b CELLD r1=900e3 r0=10000e3
xl0b16c690 l0bl16 vdd x690 x690b CELLD r1=900e3 r0=10000e3
xl0b16c691 l0bl16 vdd x691 x691b CELLD r1=900e3 r0=10000e3
xl0b16c692 l0bl16 vdd x692 x692b CELLD r1=900e3 r0=10000e3
xl0b16c693 l0bl16 vdd x693 x693b CELLD r1=900e3 r0=10000e3
xl0b16c694 l0bl16 vdd x694 x694b CELLD r1=900e3 r0=10000e3
xl0b16c695 l0bl16 vdd x695 x695b CELLD r1=900e3 r0=10000e3
xl0b16c696 l0bl16 vdd x696 x696b CELLD r1=900e3 r0=10000e3
xl0b16c697 l0bl16 vdd x697 x697b CELLD r1=900e3 r0=10000e3
xl0b16c698 l0bl16 vdd x698 x698b CELLD r1=900e3 r0=10000e3
xl0b16c699 l0bl16 vdd x699 x699b CELLD r1=10000e3 r0=900e3
xl0b16c700 l0bl16 vdd x700 x700b CELLD r1=10000e3 r0=900e3
xl0b16c701 l0bl16 vdd x701 x701b CELLD r1=900e3 r0=10000e3
xl0b16c702 l0bl16 vdd x702 x702b CELLD r1=10000e3 r0=900e3
xl0b16c703 l0bl16 vdd x703 x703b CELLD r1=900e3 r0=10000e3
xl0b16c704 l0bl16 vdd x704 x704b CELLD r1=10000e3 r0=900e3
xl0b16c705 l0bl16 vdd x705 x705b CELLD r1=900e3 r0=10000e3
xl0b16c706 l0bl16 vdd x706 x706b CELLD r1=900e3 r0=10000e3
xl0b16c707 l0bl16 vdd x707 x707b CELLD r1=900e3 r0=10000e3
xl0b16c708 l0bl16 vdd x708 x708b CELLD r1=900e3 r0=10000e3
xl0b16c709 l0bl16 vdd x709 x709b CELLD r1=900e3 r0=10000e3
xl0b16c710 l0bl16 vdd x710 x710b CELLD r1=900e3 r0=10000e3
xl0b16c711 l0bl16 vdd x711 x711b CELLD r1=900e3 r0=10000e3
xl0b16c712 l0bl16 vdd x712 x712b CELLD r1=900e3 r0=10000e3
xl0b16c713 l0bl16 vdd x713 x713b CELLD r1=900e3 r0=10000e3
xl0b16c714 l0bl16 vdd x714 x714b CELLD r1=900e3 r0=10000e3
xl0b16c715 l0bl16 vdd x715 x715b CELLD r1=900e3 r0=10000e3
xl0b16c716 l0bl16 vdd x716 x716b CELLD r1=900e3 r0=10000e3
xl0b16c717 l0bl16 vdd x717 x717b CELLD r1=900e3 r0=10000e3
xl0b16c718 l0bl16 vdd x718 x718b CELLD r1=900e3 r0=10000e3
xl0b16c719 l0bl16 vdd x719 x719b CELLD r1=10000e3 r0=900e3
xl0b16c720 l0bl16 vdd x720 x720b CELLD r1=900e3 r0=10000e3
xl0b16c721 l0bl16 vdd x721 x721b CELLD r1=900e3 r0=10000e3
xl0b16c722 l0bl16 vdd x722 x722b CELLD r1=900e3 r0=10000e3
xl0b16c723 l0bl16 vdd x723 x723b CELLD r1=10000e3 r0=900e3
xl0b16c724 l0bl16 vdd x724 x724b CELLD r1=900e3 r0=10000e3
xl0b16c725 l0bl16 vdd x725 x725b CELLD r1=10000e3 r0=900e3
xl0b16c726 l0bl16 vdd x726 x726b CELLD r1=900e3 r0=10000e3
xl0b16c727 l0bl16 vdd x727 x727b CELLD r1=900e3 r0=10000e3
xl0b16c728 l0bl16 vdd x728 x728b CELLD r1=900e3 r0=10000e3
xl0b16c729 l0bl16 vdd x729 x729b CELLD r1=900e3 r0=10000e3
xl0b16c730 l0bl16 vdd x730 x730b CELLD r1=10000e3 r0=900e3
xl0b16c731 l0bl16 vdd x731 x731b CELLD r1=10000e3 r0=900e3
xl0b16c732 l0bl16 vdd x732 x732b CELLD r1=900e3 r0=10000e3
xl0b16c733 l0bl16 vdd x733 x733b CELLD r1=900e3 r0=10000e3
xl0b16c734 l0bl16 vdd x734 x734b CELLD r1=900e3 r0=10000e3
xl0b16c735 l0bl16 vdd x735 x735b CELLD r1=900e3 r0=10000e3
xl0b16c736 l0bl16 vdd x736 x736b CELLD r1=900e3 r0=10000e3
xl0b16c737 l0bl16 vdd x737 x737b CELLD r1=900e3 r0=10000e3
xl0b16c738 l0bl16 vdd x738 x738b CELLD r1=900e3 r0=10000e3
xl0b16c739 l0bl16 vdd x739 x739b CELLD r1=10000e3 r0=900e3
xl0b16c740 l0bl16 vdd x740 x740b CELLD r1=900e3 r0=10000e3
xl0b16c741 l0bl16 vdd x741 x741b CELLD r1=900e3 r0=10000e3
xl0b16c742 l0bl16 vdd x742 x742b CELLD r1=900e3 r0=10000e3
xl0b16c743 l0bl16 vdd x743 x743b CELLD r1=900e3 r0=10000e3
xl0b16c744 l0bl16 vdd x744 x744b CELLD r1=900e3 r0=10000e3
xl0b16c745 l0bl16 vdd x745 x745b CELLD r1=900e3 r0=10000e3
xl0b16c746 l0bl16 vdd x746 x746b CELLD r1=10000e3 r0=900e3
xl0b16c747 l0bl16 vdd x747 x747b CELLD r1=10000e3 r0=900e3
xl0b16c748 l0bl16 vdd x748 x748b CELLD r1=900e3 r0=10000e3
xl0b16c749 l0bl16 vdd x749 x749b CELLD r1=900e3 r0=10000e3
xl0b16c750 l0bl16 vdd x750 x750b CELLD r1=900e3 r0=10000e3
xl0b16c751 l0bl16 vdd x751 x751b CELLD r1=900e3 r0=10000e3
xl0b16c752 l0bl16 vdd x752 x752b CELLD r1=10000e3 r0=900e3
xl0b16c753 l0bl16 vdd x753 x753b CELLD r1=10000e3 r0=900e3
xl0b16c754 l0bl16 vdd x754 x754b CELLD r1=900e3 r0=10000e3
xl0b16c755 l0bl16 vdd x755 x755b CELLD r1=10000e3 r0=900e3
xl0b16c756 l0bl16 vdd x756 x756b CELLD r1=10000e3 r0=900e3
xl0b16c757 l0bl16 vdd x757 x757b CELLD r1=900e3 r0=10000e3
xl0b16c758 l0bl16 vdd x758 x758b CELLD r1=900e3 r0=10000e3
xl0b16c759 l0bl16 vdd x759 x759b CELLD r1=10000e3 r0=900e3
xl0b16c760 l0bl16 vdd x760 x760b CELLD r1=10000e3 r0=900e3
xl0b16c761 l0bl16 vdd x761 x761b CELLD r1=10000e3 r0=900e3
xl0b16c762 l0bl16 vdd x762 x762b CELLD r1=10000e3 r0=900e3
xl0b16c763 l0bl16 vdd x763 x763b CELLD r1=900e3 r0=10000e3
xl0b16c764 l0bl16 vdd x764 x764b CELLD r1=900e3 r0=10000e3
xl0b16c765 l0bl16 vdd x765 x765b CELLD r1=900e3 r0=10000e3
xl0b16c766 l0bl16 vdd x766 x766b CELLD r1=10000e3 r0=900e3
xl0b16c767 l0bl16 vdd x767 x767b CELLD r1=900e3 r0=10000e3
xl0b16c768 l0bl16 vdd x768 x768b CELLD r1=900e3 r0=10000e3
xl0b16c769 l0bl16 vdd x769 x769b CELLD r1=10000e3 r0=900e3
xl0b16c770 l0bl16 vdd x770 x770b CELLD r1=10000e3 r0=900e3
xl0b16c771 l0bl16 vdd x771 x771b CELLD r1=900e3 r0=10000e3
xl0b16c772 l0bl16 vdd x772 x772b CELLD r1=900e3 r0=10000e3
xl0b16c773 l0bl16 vdd x773 x773b CELLD r1=900e3 r0=10000e3
xl0b16c774 l0bl16 vdd x774 x774b CELLD r1=900e3 r0=10000e3
xl0b16c775 l0bl16 vdd x775 x775b CELLD r1=900e3 r0=10000e3
xl0b16c776 l0bl16 vdd x776 x776b CELLD r1=900e3 r0=10000e3
xl0b16c777 l0bl16 vdd x777 x777b CELLD r1=10000e3 r0=900e3
xl0b16c778 l0bl16 vdd x778 x778b CELLD r1=10000e3 r0=900e3
xl0b16c779 l0bl16 vdd x779 x779b CELLD r1=10000e3 r0=900e3
xl0b16c780 l0bl16 vdd x780 x780b CELLD r1=10000e3 r0=900e3
xl0b16c781 l0bl16 vdd x781 x781b CELLD r1=900e3 r0=10000e3
xl0b16c782 l0bl16 vdd x782 x782b CELLD r1=900e3 r0=10000e3
xl0b16c783 l0bl16 vdd x783 x783b CELLD r1=10000e3 r0=900e3
xl0b17c0 l0bl17 vdd x0 x0b CELLD r1=900e3 r0=10000e3
xl0b17c1 l0bl17 vdd x1 x1b CELLD r1=900e3 r0=10000e3
xl0b17c2 l0bl17 vdd x2 x2b CELLD r1=900e3 r0=10000e3
xl0b17c3 l0bl17 vdd x3 x3b CELLD r1=900e3 r0=10000e3
xl0b17c4 l0bl17 vdd x4 x4b CELLD r1=10000e3 r0=900e3
xl0b17c5 l0bl17 vdd x5 x5b CELLD r1=900e3 r0=10000e3
xl0b17c6 l0bl17 vdd x6 x6b CELLD r1=900e3 r0=10000e3
xl0b17c7 l0bl17 vdd x7 x7b CELLD r1=10000e3 r0=900e3
xl0b17c8 l0bl17 vdd x8 x8b CELLD r1=10000e3 r0=900e3
xl0b17c9 l0bl17 vdd x9 x9b CELLD r1=900e3 r0=10000e3
xl0b17c10 l0bl17 vdd x10 x10b CELLD r1=900e3 r0=10000e3
xl0b17c11 l0bl17 vdd x11 x11b CELLD r1=900e3 r0=10000e3
xl0b17c12 l0bl17 vdd x12 x12b CELLD r1=900e3 r0=10000e3
xl0b17c13 l0bl17 vdd x13 x13b CELLD r1=900e3 r0=10000e3
xl0b17c14 l0bl17 vdd x14 x14b CELLD r1=900e3 r0=10000e3
xl0b17c15 l0bl17 vdd x15 x15b CELLD r1=900e3 r0=10000e3
xl0b17c16 l0bl17 vdd x16 x16b CELLD r1=900e3 r0=10000e3
xl0b17c17 l0bl17 vdd x17 x17b CELLD r1=900e3 r0=10000e3
xl0b17c18 l0bl17 vdd x18 x18b CELLD r1=900e3 r0=10000e3
xl0b17c19 l0bl17 vdd x19 x19b CELLD r1=900e3 r0=10000e3
xl0b17c20 l0bl17 vdd x20 x20b CELLD r1=10000e3 r0=900e3
xl0b17c21 l0bl17 vdd x21 x21b CELLD r1=900e3 r0=10000e3
xl0b17c22 l0bl17 vdd x22 x22b CELLD r1=900e3 r0=10000e3
xl0b17c23 l0bl17 vdd x23 x23b CELLD r1=900e3 r0=10000e3
xl0b17c24 l0bl17 vdd x24 x24b CELLD r1=10000e3 r0=900e3
xl0b17c25 l0bl17 vdd x25 x25b CELLD r1=900e3 r0=10000e3
xl0b17c26 l0bl17 vdd x26 x26b CELLD r1=900e3 r0=10000e3
xl0b17c27 l0bl17 vdd x27 x27b CELLD r1=10000e3 r0=900e3
xl0b17c28 l0bl17 vdd x28 x28b CELLD r1=900e3 r0=10000e3
xl0b17c29 l0bl17 vdd x29 x29b CELLD r1=900e3 r0=10000e3
xl0b17c30 l0bl17 vdd x30 x30b CELLD r1=10000e3 r0=900e3
xl0b17c31 l0bl17 vdd x31 x31b CELLD r1=900e3 r0=10000e3
xl0b17c32 l0bl17 vdd x32 x32b CELLD r1=900e3 r0=10000e3
xl0b17c33 l0bl17 vdd x33 x33b CELLD r1=900e3 r0=10000e3
xl0b17c34 l0bl17 vdd x34 x34b CELLD r1=900e3 r0=10000e3
xl0b17c35 l0bl17 vdd x35 x35b CELLD r1=900e3 r0=10000e3
xl0b17c36 l0bl17 vdd x36 x36b CELLD r1=900e3 r0=10000e3
xl0b17c37 l0bl17 vdd x37 x37b CELLD r1=10000e3 r0=900e3
xl0b17c38 l0bl17 vdd x38 x38b CELLD r1=900e3 r0=10000e3
xl0b17c39 l0bl17 vdd x39 x39b CELLD r1=900e3 r0=10000e3
xl0b17c40 l0bl17 vdd x40 x40b CELLD r1=10000e3 r0=900e3
xl0b17c41 l0bl17 vdd x41 x41b CELLD r1=900e3 r0=10000e3
xl0b17c42 l0bl17 vdd x42 x42b CELLD r1=900e3 r0=10000e3
xl0b17c43 l0bl17 vdd x43 x43b CELLD r1=900e3 r0=10000e3
xl0b17c44 l0bl17 vdd x44 x44b CELLD r1=900e3 r0=10000e3
xl0b17c45 l0bl17 vdd x45 x45b CELLD r1=10000e3 r0=900e3
xl0b17c46 l0bl17 vdd x46 x46b CELLD r1=900e3 r0=10000e3
xl0b17c47 l0bl17 vdd x47 x47b CELLD r1=10000e3 r0=900e3
xl0b17c48 l0bl17 vdd x48 x48b CELLD r1=10000e3 r0=900e3
xl0b17c49 l0bl17 vdd x49 x49b CELLD r1=10000e3 r0=900e3
xl0b17c50 l0bl17 vdd x50 x50b CELLD r1=900e3 r0=10000e3
xl0b17c51 l0bl17 vdd x51 x51b CELLD r1=10000e3 r0=900e3
xl0b17c52 l0bl17 vdd x52 x52b CELLD r1=900e3 r0=10000e3
xl0b17c53 l0bl17 vdd x53 x53b CELLD r1=10000e3 r0=900e3
xl0b17c54 l0bl17 vdd x54 x54b CELLD r1=900e3 r0=10000e3
xl0b17c55 l0bl17 vdd x55 x55b CELLD r1=10000e3 r0=900e3
xl0b17c56 l0bl17 vdd x56 x56b CELLD r1=900e3 r0=10000e3
xl0b17c57 l0bl17 vdd x57 x57b CELLD r1=900e3 r0=10000e3
xl0b17c58 l0bl17 vdd x58 x58b CELLD r1=10000e3 r0=900e3
xl0b17c59 l0bl17 vdd x59 x59b CELLD r1=900e3 r0=10000e3
xl0b17c60 l0bl17 vdd x60 x60b CELLD r1=900e3 r0=10000e3
xl0b17c61 l0bl17 vdd x61 x61b CELLD r1=900e3 r0=10000e3
xl0b17c62 l0bl17 vdd x62 x62b CELLD r1=900e3 r0=10000e3
xl0b17c63 l0bl17 vdd x63 x63b CELLD r1=10000e3 r0=900e3
xl0b17c64 l0bl17 vdd x64 x64b CELLD r1=10000e3 r0=900e3
xl0b17c65 l0bl17 vdd x65 x65b CELLD r1=900e3 r0=10000e3
xl0b17c66 l0bl17 vdd x66 x66b CELLD r1=10000e3 r0=900e3
xl0b17c67 l0bl17 vdd x67 x67b CELLD r1=900e3 r0=10000e3
xl0b17c68 l0bl17 vdd x68 x68b CELLD r1=10000e3 r0=900e3
xl0b17c69 l0bl17 vdd x69 x69b CELLD r1=10000e3 r0=900e3
xl0b17c70 l0bl17 vdd x70 x70b CELLD r1=900e3 r0=10000e3
xl0b17c71 l0bl17 vdd x71 x71b CELLD r1=10000e3 r0=900e3
xl0b17c72 l0bl17 vdd x72 x72b CELLD r1=10000e3 r0=900e3
xl0b17c73 l0bl17 vdd x73 x73b CELLD r1=10000e3 r0=900e3
xl0b17c74 l0bl17 vdd x74 x74b CELLD r1=900e3 r0=10000e3
xl0b17c75 l0bl17 vdd x75 x75b CELLD r1=900e3 r0=10000e3
xl0b17c76 l0bl17 vdd x76 x76b CELLD r1=900e3 r0=10000e3
xl0b17c77 l0bl17 vdd x77 x77b CELLD r1=900e3 r0=10000e3
xl0b17c78 l0bl17 vdd x78 x78b CELLD r1=900e3 r0=10000e3
xl0b17c79 l0bl17 vdd x79 x79b CELLD r1=900e3 r0=10000e3
xl0b17c80 l0bl17 vdd x80 x80b CELLD r1=900e3 r0=10000e3
xl0b17c81 l0bl17 vdd x81 x81b CELLD r1=900e3 r0=10000e3
xl0b17c82 l0bl17 vdd x82 x82b CELLD r1=900e3 r0=10000e3
xl0b17c83 l0bl17 vdd x83 x83b CELLD r1=10000e3 r0=900e3
xl0b17c84 l0bl17 vdd x84 x84b CELLD r1=10000e3 r0=900e3
xl0b17c85 l0bl17 vdd x85 x85b CELLD r1=900e3 r0=10000e3
xl0b17c86 l0bl17 vdd x86 x86b CELLD r1=10000e3 r0=900e3
xl0b17c87 l0bl17 vdd x87 x87b CELLD r1=900e3 r0=10000e3
xl0b17c88 l0bl17 vdd x88 x88b CELLD r1=900e3 r0=10000e3
xl0b17c89 l0bl17 vdd x89 x89b CELLD r1=10000e3 r0=900e3
xl0b17c90 l0bl17 vdd x90 x90b CELLD r1=900e3 r0=10000e3
xl0b17c91 l0bl17 vdd x91 x91b CELLD r1=10000e3 r0=900e3
xl0b17c92 l0bl17 vdd x92 x92b CELLD r1=10000e3 r0=900e3
xl0b17c93 l0bl17 vdd x93 x93b CELLD r1=10000e3 r0=900e3
xl0b17c94 l0bl17 vdd x94 x94b CELLD r1=10000e3 r0=900e3
xl0b17c95 l0bl17 vdd x95 x95b CELLD r1=10000e3 r0=900e3
xl0b17c96 l0bl17 vdd x96 x96b CELLD r1=10000e3 r0=900e3
xl0b17c97 l0bl17 vdd x97 x97b CELLD r1=10000e3 r0=900e3
xl0b17c98 l0bl17 vdd x98 x98b CELLD r1=10000e3 r0=900e3
xl0b17c99 l0bl17 vdd x99 x99b CELLD r1=10000e3 r0=900e3
xl0b17c100 l0bl17 vdd x100 x100b CELLD r1=10000e3 r0=900e3
xl0b17c101 l0bl17 vdd x101 x101b CELLD r1=10000e3 r0=900e3
xl0b17c102 l0bl17 vdd x102 x102b CELLD r1=900e3 r0=10000e3
xl0b17c103 l0bl17 vdd x103 x103b CELLD r1=900e3 r0=10000e3
xl0b17c104 l0bl17 vdd x104 x104b CELLD r1=10000e3 r0=900e3
xl0b17c105 l0bl17 vdd x105 x105b CELLD r1=900e3 r0=10000e3
xl0b17c106 l0bl17 vdd x106 x106b CELLD r1=900e3 r0=10000e3
xl0b17c107 l0bl17 vdd x107 x107b CELLD r1=900e3 r0=10000e3
xl0b17c108 l0bl17 vdd x108 x108b CELLD r1=900e3 r0=10000e3
xl0b17c109 l0bl17 vdd x109 x109b CELLD r1=900e3 r0=10000e3
xl0b17c110 l0bl17 vdd x110 x110b CELLD r1=900e3 r0=10000e3
xl0b17c111 l0bl17 vdd x111 x111b CELLD r1=900e3 r0=10000e3
xl0b17c112 l0bl17 vdd x112 x112b CELLD r1=900e3 r0=10000e3
xl0b17c113 l0bl17 vdd x113 x113b CELLD r1=10000e3 r0=900e3
xl0b17c114 l0bl17 vdd x114 x114b CELLD r1=900e3 r0=10000e3
xl0b17c115 l0bl17 vdd x115 x115b CELLD r1=10000e3 r0=900e3
xl0b17c116 l0bl17 vdd x116 x116b CELLD r1=900e3 r0=10000e3
xl0b17c117 l0bl17 vdd x117 x117b CELLD r1=10000e3 r0=900e3
xl0b17c118 l0bl17 vdd x118 x118b CELLD r1=900e3 r0=10000e3
xl0b17c119 l0bl17 vdd x119 x119b CELLD r1=900e3 r0=10000e3
xl0b17c120 l0bl17 vdd x120 x120b CELLD r1=10000e3 r0=900e3
xl0b17c121 l0bl17 vdd x121 x121b CELLD r1=10000e3 r0=900e3
xl0b17c122 l0bl17 vdd x122 x122b CELLD r1=10000e3 r0=900e3
xl0b17c123 l0bl17 vdd x123 x123b CELLD r1=10000e3 r0=900e3
xl0b17c124 l0bl17 vdd x124 x124b CELLD r1=10000e3 r0=900e3
xl0b17c125 l0bl17 vdd x125 x125b CELLD r1=10000e3 r0=900e3
xl0b17c126 l0bl17 vdd x126 x126b CELLD r1=10000e3 r0=900e3
xl0b17c127 l0bl17 vdd x127 x127b CELLD r1=10000e3 r0=900e3
xl0b17c128 l0bl17 vdd x128 x128b CELLD r1=10000e3 r0=900e3
xl0b17c129 l0bl17 vdd x129 x129b CELLD r1=10000e3 r0=900e3
xl0b17c130 l0bl17 vdd x130 x130b CELLD r1=10000e3 r0=900e3
xl0b17c131 l0bl17 vdd x131 x131b CELLD r1=900e3 r0=10000e3
xl0b17c132 l0bl17 vdd x132 x132b CELLD r1=900e3 r0=10000e3
xl0b17c133 l0bl17 vdd x133 x133b CELLD r1=900e3 r0=10000e3
xl0b17c134 l0bl17 vdd x134 x134b CELLD r1=900e3 r0=10000e3
xl0b17c135 l0bl17 vdd x135 x135b CELLD r1=10000e3 r0=900e3
xl0b17c136 l0bl17 vdd x136 x136b CELLD r1=10000e3 r0=900e3
xl0b17c137 l0bl17 vdd x137 x137b CELLD r1=900e3 r0=10000e3
xl0b17c138 l0bl17 vdd x138 x138b CELLD r1=900e3 r0=10000e3
xl0b17c139 l0bl17 vdd x139 x139b CELLD r1=10000e3 r0=900e3
xl0b17c140 l0bl17 vdd x140 x140b CELLD r1=10000e3 r0=900e3
xl0b17c141 l0bl17 vdd x141 x141b CELLD r1=900e3 r0=10000e3
xl0b17c142 l0bl17 vdd x142 x142b CELLD r1=10000e3 r0=900e3
xl0b17c143 l0bl17 vdd x143 x143b CELLD r1=900e3 r0=10000e3
xl0b17c144 l0bl17 vdd x144 x144b CELLD r1=10000e3 r0=900e3
xl0b17c145 l0bl17 vdd x145 x145b CELLD r1=10000e3 r0=900e3
xl0b17c146 l0bl17 vdd x146 x146b CELLD r1=10000e3 r0=900e3
xl0b17c147 l0bl17 vdd x147 x147b CELLD r1=10000e3 r0=900e3
xl0b17c148 l0bl17 vdd x148 x148b CELLD r1=10000e3 r0=900e3
xl0b17c149 l0bl17 vdd x149 x149b CELLD r1=10000e3 r0=900e3
xl0b17c150 l0bl17 vdd x150 x150b CELLD r1=10000e3 r0=900e3
xl0b17c151 l0bl17 vdd x151 x151b CELLD r1=10000e3 r0=900e3
xl0b17c152 l0bl17 vdd x152 x152b CELLD r1=10000e3 r0=900e3
xl0b17c153 l0bl17 vdd x153 x153b CELLD r1=10000e3 r0=900e3
xl0b17c154 l0bl17 vdd x154 x154b CELLD r1=900e3 r0=10000e3
xl0b17c155 l0bl17 vdd x155 x155b CELLD r1=10000e3 r0=900e3
xl0b17c156 l0bl17 vdd x156 x156b CELLD r1=10000e3 r0=900e3
xl0b17c157 l0bl17 vdd x157 x157b CELLD r1=10000e3 r0=900e3
xl0b17c158 l0bl17 vdd x158 x158b CELLD r1=900e3 r0=10000e3
xl0b17c159 l0bl17 vdd x159 x159b CELLD r1=900e3 r0=10000e3
xl0b17c160 l0bl17 vdd x160 x160b CELLD r1=900e3 r0=10000e3
xl0b17c161 l0bl17 vdd x161 x161b CELLD r1=900e3 r0=10000e3
xl0b17c162 l0bl17 vdd x162 x162b CELLD r1=900e3 r0=10000e3
xl0b17c163 l0bl17 vdd x163 x163b CELLD r1=900e3 r0=10000e3
xl0b17c164 l0bl17 vdd x164 x164b CELLD r1=900e3 r0=10000e3
xl0b17c165 l0bl17 vdd x165 x165b CELLD r1=900e3 r0=10000e3
xl0b17c166 l0bl17 vdd x166 x166b CELLD r1=900e3 r0=10000e3
xl0b17c167 l0bl17 vdd x167 x167b CELLD r1=900e3 r0=10000e3
xl0b17c168 l0bl17 vdd x168 x168b CELLD r1=10000e3 r0=900e3
xl0b17c169 l0bl17 vdd x169 x169b CELLD r1=900e3 r0=10000e3
xl0b17c170 l0bl17 vdd x170 x170b CELLD r1=900e3 r0=10000e3
xl0b17c171 l0bl17 vdd x171 x171b CELLD r1=900e3 r0=10000e3
xl0b17c172 l0bl17 vdd x172 x172b CELLD r1=900e3 r0=10000e3
xl0b17c173 l0bl17 vdd x173 x173b CELLD r1=900e3 r0=10000e3
xl0b17c174 l0bl17 vdd x174 x174b CELLD r1=900e3 r0=10000e3
xl0b17c175 l0bl17 vdd x175 x175b CELLD r1=10000e3 r0=900e3
xl0b17c176 l0bl17 vdd x176 x176b CELLD r1=10000e3 r0=900e3
xl0b17c177 l0bl17 vdd x177 x177b CELLD r1=10000e3 r0=900e3
xl0b17c178 l0bl17 vdd x178 x178b CELLD r1=10000e3 r0=900e3
xl0b17c179 l0bl17 vdd x179 x179b CELLD r1=10000e3 r0=900e3
xl0b17c180 l0bl17 vdd x180 x180b CELLD r1=10000e3 r0=900e3
xl0b17c181 l0bl17 vdd x181 x181b CELLD r1=900e3 r0=10000e3
xl0b17c182 l0bl17 vdd x182 x182b CELLD r1=10000e3 r0=900e3
xl0b17c183 l0bl17 vdd x183 x183b CELLD r1=10000e3 r0=900e3
xl0b17c184 l0bl17 vdd x184 x184b CELLD r1=10000e3 r0=900e3
xl0b17c185 l0bl17 vdd x185 x185b CELLD r1=900e3 r0=10000e3
xl0b17c186 l0bl17 vdd x186 x186b CELLD r1=900e3 r0=10000e3
xl0b17c187 l0bl17 vdd x187 x187b CELLD r1=900e3 r0=10000e3
xl0b17c188 l0bl17 vdd x188 x188b CELLD r1=900e3 r0=10000e3
xl0b17c189 l0bl17 vdd x189 x189b CELLD r1=900e3 r0=10000e3
xl0b17c190 l0bl17 vdd x190 x190b CELLD r1=900e3 r0=10000e3
xl0b17c191 l0bl17 vdd x191 x191b CELLD r1=900e3 r0=10000e3
xl0b17c192 l0bl17 vdd x192 x192b CELLD r1=900e3 r0=10000e3
xl0b17c193 l0bl17 vdd x193 x193b CELLD r1=10000e3 r0=900e3
xl0b17c194 l0bl17 vdd x194 x194b CELLD r1=900e3 r0=10000e3
xl0b17c195 l0bl17 vdd x195 x195b CELLD r1=900e3 r0=10000e3
xl0b17c196 l0bl17 vdd x196 x196b CELLD r1=900e3 r0=10000e3
xl0b17c197 l0bl17 vdd x197 x197b CELLD r1=900e3 r0=10000e3
xl0b17c198 l0bl17 vdd x198 x198b CELLD r1=10000e3 r0=900e3
xl0b17c199 l0bl17 vdd x199 x199b CELLD r1=900e3 r0=10000e3
xl0b17c200 l0bl17 vdd x200 x200b CELLD r1=900e3 r0=10000e3
xl0b17c201 l0bl17 vdd x201 x201b CELLD r1=900e3 r0=10000e3
xl0b17c202 l0bl17 vdd x202 x202b CELLD r1=10000e3 r0=900e3
xl0b17c203 l0bl17 vdd x203 x203b CELLD r1=10000e3 r0=900e3
xl0b17c204 l0bl17 vdd x204 x204b CELLD r1=10000e3 r0=900e3
xl0b17c205 l0bl17 vdd x205 x205b CELLD r1=10000e3 r0=900e3
xl0b17c206 l0bl17 vdd x206 x206b CELLD r1=10000e3 r0=900e3
xl0b17c207 l0bl17 vdd x207 x207b CELLD r1=10000e3 r0=900e3
xl0b17c208 l0bl17 vdd x208 x208b CELLD r1=10000e3 r0=900e3
xl0b17c209 l0bl17 vdd x209 x209b CELLD r1=10000e3 r0=900e3
xl0b17c210 l0bl17 vdd x210 x210b CELLD r1=10000e3 r0=900e3
xl0b17c211 l0bl17 vdd x211 x211b CELLD r1=10000e3 r0=900e3
xl0b17c212 l0bl17 vdd x212 x212b CELLD r1=900e3 r0=10000e3
xl0b17c213 l0bl17 vdd x213 x213b CELLD r1=900e3 r0=10000e3
xl0b17c214 l0bl17 vdd x214 x214b CELLD r1=900e3 r0=10000e3
xl0b17c215 l0bl17 vdd x215 x215b CELLD r1=10000e3 r0=900e3
xl0b17c216 l0bl17 vdd x216 x216b CELLD r1=10000e3 r0=900e3
xl0b17c217 l0bl17 vdd x217 x217b CELLD r1=10000e3 r0=900e3
xl0b17c218 l0bl17 vdd x218 x218b CELLD r1=10000e3 r0=900e3
xl0b17c219 l0bl17 vdd x219 x219b CELLD r1=900e3 r0=10000e3
xl0b17c220 l0bl17 vdd x220 x220b CELLD r1=10000e3 r0=900e3
xl0b17c221 l0bl17 vdd x221 x221b CELLD r1=10000e3 r0=900e3
xl0b17c222 l0bl17 vdd x222 x222b CELLD r1=900e3 r0=10000e3
xl0b17c223 l0bl17 vdd x223 x223b CELLD r1=10000e3 r0=900e3
xl0b17c224 l0bl17 vdd x224 x224b CELLD r1=10000e3 r0=900e3
xl0b17c225 l0bl17 vdd x225 x225b CELLD r1=10000e3 r0=900e3
xl0b17c226 l0bl17 vdd x226 x226b CELLD r1=10000e3 r0=900e3
xl0b17c227 l0bl17 vdd x227 x227b CELLD r1=900e3 r0=10000e3
xl0b17c228 l0bl17 vdd x228 x228b CELLD r1=10000e3 r0=900e3
xl0b17c229 l0bl17 vdd x229 x229b CELLD r1=900e3 r0=10000e3
xl0b17c230 l0bl17 vdd x230 x230b CELLD r1=10000e3 r0=900e3
xl0b17c231 l0bl17 vdd x231 x231b CELLD r1=10000e3 r0=900e3
xl0b17c232 l0bl17 vdd x232 x232b CELLD r1=10000e3 r0=900e3
xl0b17c233 l0bl17 vdd x233 x233b CELLD r1=10000e3 r0=900e3
xl0b17c234 l0bl17 vdd x234 x234b CELLD r1=10000e3 r0=900e3
xl0b17c235 l0bl17 vdd x235 x235b CELLD r1=10000e3 r0=900e3
xl0b17c236 l0bl17 vdd x236 x236b CELLD r1=10000e3 r0=900e3
xl0b17c237 l0bl17 vdd x237 x237b CELLD r1=10000e3 r0=900e3
xl0b17c238 l0bl17 vdd x238 x238b CELLD r1=900e3 r0=10000e3
xl0b17c239 l0bl17 vdd x239 x239b CELLD r1=900e3 r0=10000e3
xl0b17c240 l0bl17 vdd x240 x240b CELLD r1=900e3 r0=10000e3
xl0b17c241 l0bl17 vdd x241 x241b CELLD r1=900e3 r0=10000e3
xl0b17c242 l0bl17 vdd x242 x242b CELLD r1=900e3 r0=10000e3
xl0b17c243 l0bl17 vdd x243 x243b CELLD r1=10000e3 r0=900e3
xl0b17c244 l0bl17 vdd x244 x244b CELLD r1=10000e3 r0=900e3
xl0b17c245 l0bl17 vdd x245 x245b CELLD r1=10000e3 r0=900e3
xl0b17c246 l0bl17 vdd x246 x246b CELLD r1=10000e3 r0=900e3
xl0b17c247 l0bl17 vdd x247 x247b CELLD r1=10000e3 r0=900e3
xl0b17c248 l0bl17 vdd x248 x248b CELLD r1=10000e3 r0=900e3
xl0b17c249 l0bl17 vdd x249 x249b CELLD r1=10000e3 r0=900e3
xl0b17c250 l0bl17 vdd x250 x250b CELLD r1=10000e3 r0=900e3
xl0b17c251 l0bl17 vdd x251 x251b CELLD r1=10000e3 r0=900e3
xl0b17c252 l0bl17 vdd x252 x252b CELLD r1=10000e3 r0=900e3
xl0b17c253 l0bl17 vdd x253 x253b CELLD r1=900e3 r0=10000e3
xl0b17c254 l0bl17 vdd x254 x254b CELLD r1=10000e3 r0=900e3
xl0b17c255 l0bl17 vdd x255 x255b CELLD r1=10000e3 r0=900e3
xl0b17c256 l0bl17 vdd x256 x256b CELLD r1=900e3 r0=10000e3
xl0b17c257 l0bl17 vdd x257 x257b CELLD r1=10000e3 r0=900e3
xl0b17c258 l0bl17 vdd x258 x258b CELLD r1=10000e3 r0=900e3
xl0b17c259 l0bl17 vdd x259 x259b CELLD r1=10000e3 r0=900e3
xl0b17c260 l0bl17 vdd x260 x260b CELLD r1=10000e3 r0=900e3
xl0b17c261 l0bl17 vdd x261 x261b CELLD r1=10000e3 r0=900e3
xl0b17c262 l0bl17 vdd x262 x262b CELLD r1=10000e3 r0=900e3
xl0b17c263 l0bl17 vdd x263 x263b CELLD r1=900e3 r0=10000e3
xl0b17c264 l0bl17 vdd x264 x264b CELLD r1=900e3 r0=10000e3
xl0b17c265 l0bl17 vdd x265 x265b CELLD r1=900e3 r0=10000e3
xl0b17c266 l0bl17 vdd x266 x266b CELLD r1=10000e3 r0=900e3
xl0b17c267 l0bl17 vdd x267 x267b CELLD r1=10000e3 r0=900e3
xl0b17c268 l0bl17 vdd x268 x268b CELLD r1=10000e3 r0=900e3
xl0b17c269 l0bl17 vdd x269 x269b CELLD r1=10000e3 r0=900e3
xl0b17c270 l0bl17 vdd x270 x270b CELLD r1=10000e3 r0=900e3
xl0b17c271 l0bl17 vdd x271 x271b CELLD r1=10000e3 r0=900e3
xl0b17c272 l0bl17 vdd x272 x272b CELLD r1=10000e3 r0=900e3
xl0b17c273 l0bl17 vdd x273 x273b CELLD r1=10000e3 r0=900e3
xl0b17c274 l0bl17 vdd x274 x274b CELLD r1=10000e3 r0=900e3
xl0b17c275 l0bl17 vdd x275 x275b CELLD r1=10000e3 r0=900e3
xl0b17c276 l0bl17 vdd x276 x276b CELLD r1=10000e3 r0=900e3
xl0b17c277 l0bl17 vdd x277 x277b CELLD r1=10000e3 r0=900e3
xl0b17c278 l0bl17 vdd x278 x278b CELLD r1=10000e3 r0=900e3
xl0b17c279 l0bl17 vdd x279 x279b CELLD r1=900e3 r0=10000e3
xl0b17c280 l0bl17 vdd x280 x280b CELLD r1=900e3 r0=10000e3
xl0b17c281 l0bl17 vdd x281 x281b CELLD r1=10000e3 r0=900e3
xl0b17c282 l0bl17 vdd x282 x282b CELLD r1=10000e3 r0=900e3
xl0b17c283 l0bl17 vdd x283 x283b CELLD r1=900e3 r0=10000e3
xl0b17c284 l0bl17 vdd x284 x284b CELLD r1=10000e3 r0=900e3
xl0b17c285 l0bl17 vdd x285 x285b CELLD r1=10000e3 r0=900e3
xl0b17c286 l0bl17 vdd x286 x286b CELLD r1=10000e3 r0=900e3
xl0b17c287 l0bl17 vdd x287 x287b CELLD r1=10000e3 r0=900e3
xl0b17c288 l0bl17 vdd x288 x288b CELLD r1=10000e3 r0=900e3
xl0b17c289 l0bl17 vdd x289 x289b CELLD r1=10000e3 r0=900e3
xl0b17c290 l0bl17 vdd x290 x290b CELLD r1=900e3 r0=10000e3
xl0b17c291 l0bl17 vdd x291 x291b CELLD r1=900e3 r0=10000e3
xl0b17c292 l0bl17 vdd x292 x292b CELLD r1=900e3 r0=10000e3
xl0b17c293 l0bl17 vdd x293 x293b CELLD r1=900e3 r0=10000e3
xl0b17c294 l0bl17 vdd x294 x294b CELLD r1=900e3 r0=10000e3
xl0b17c295 l0bl17 vdd x295 x295b CELLD r1=900e3 r0=10000e3
xl0b17c296 l0bl17 vdd x296 x296b CELLD r1=10000e3 r0=900e3
xl0b17c297 l0bl17 vdd x297 x297b CELLD r1=10000e3 r0=900e3
xl0b17c298 l0bl17 vdd x298 x298b CELLD r1=10000e3 r0=900e3
xl0b17c299 l0bl17 vdd x299 x299b CELLD r1=10000e3 r0=900e3
xl0b17c300 l0bl17 vdd x300 x300b CELLD r1=10000e3 r0=900e3
xl0b17c301 l0bl17 vdd x301 x301b CELLD r1=10000e3 r0=900e3
xl0b17c302 l0bl17 vdd x302 x302b CELLD r1=10000e3 r0=900e3
xl0b17c303 l0bl17 vdd x303 x303b CELLD r1=10000e3 r0=900e3
xl0b17c304 l0bl17 vdd x304 x304b CELLD r1=10000e3 r0=900e3
xl0b17c305 l0bl17 vdd x305 x305b CELLD r1=10000e3 r0=900e3
xl0b17c306 l0bl17 vdd x306 x306b CELLD r1=900e3 r0=10000e3
xl0b17c307 l0bl17 vdd x307 x307b CELLD r1=10000e3 r0=900e3
xl0b17c308 l0bl17 vdd x308 x308b CELLD r1=900e3 r0=10000e3
xl0b17c309 l0bl17 vdd x309 x309b CELLD r1=900e3 r0=10000e3
xl0b17c310 l0bl17 vdd x310 x310b CELLD r1=10000e3 r0=900e3
xl0b17c311 l0bl17 vdd x311 x311b CELLD r1=10000e3 r0=900e3
xl0b17c312 l0bl17 vdd x312 x312b CELLD r1=10000e3 r0=900e3
xl0b17c313 l0bl17 vdd x313 x313b CELLD r1=10000e3 r0=900e3
xl0b17c314 l0bl17 vdd x314 x314b CELLD r1=10000e3 r0=900e3
xl0b17c315 l0bl17 vdd x315 x315b CELLD r1=10000e3 r0=900e3
xl0b17c316 l0bl17 vdd x316 x316b CELLD r1=10000e3 r0=900e3
xl0b17c317 l0bl17 vdd x317 x317b CELLD r1=900e3 r0=10000e3
xl0b17c318 l0bl17 vdd x318 x318b CELLD r1=900e3 r0=10000e3
xl0b17c319 l0bl17 vdd x319 x319b CELLD r1=900e3 r0=10000e3
xl0b17c320 l0bl17 vdd x320 x320b CELLD r1=900e3 r0=10000e3
xl0b17c321 l0bl17 vdd x321 x321b CELLD r1=900e3 r0=10000e3
xl0b17c322 l0bl17 vdd x322 x322b CELLD r1=900e3 r0=10000e3
xl0b17c323 l0bl17 vdd x323 x323b CELLD r1=900e3 r0=10000e3
xl0b17c324 l0bl17 vdd x324 x324b CELLD r1=900e3 r0=10000e3
xl0b17c325 l0bl17 vdd x325 x325b CELLD r1=900e3 r0=10000e3
xl0b17c326 l0bl17 vdd x326 x326b CELLD r1=10000e3 r0=900e3
xl0b17c327 l0bl17 vdd x327 x327b CELLD r1=10000e3 r0=900e3
xl0b17c328 l0bl17 vdd x328 x328b CELLD r1=10000e3 r0=900e3
xl0b17c329 l0bl17 vdd x329 x329b CELLD r1=10000e3 r0=900e3
xl0b17c330 l0bl17 vdd x330 x330b CELLD r1=10000e3 r0=900e3
xl0b17c331 l0bl17 vdd x331 x331b CELLD r1=10000e3 r0=900e3
xl0b17c332 l0bl17 vdd x332 x332b CELLD r1=10000e3 r0=900e3
xl0b17c333 l0bl17 vdd x333 x333b CELLD r1=10000e3 r0=900e3
xl0b17c334 l0bl17 vdd x334 x334b CELLD r1=900e3 r0=10000e3
xl0b17c335 l0bl17 vdd x335 x335b CELLD r1=900e3 r0=10000e3
xl0b17c336 l0bl17 vdd x336 x336b CELLD r1=10000e3 r0=900e3
xl0b17c337 l0bl17 vdd x337 x337b CELLD r1=900e3 r0=10000e3
xl0b17c338 l0bl17 vdd x338 x338b CELLD r1=10000e3 r0=900e3
xl0b17c339 l0bl17 vdd x339 x339b CELLD r1=10000e3 r0=900e3
xl0b17c340 l0bl17 vdd x340 x340b CELLD r1=10000e3 r0=900e3
xl0b17c341 l0bl17 vdd x341 x341b CELLD r1=10000e3 r0=900e3
xl0b17c342 l0bl17 vdd x342 x342b CELLD r1=10000e3 r0=900e3
xl0b17c343 l0bl17 vdd x343 x343b CELLD r1=10000e3 r0=900e3
xl0b17c344 l0bl17 vdd x344 x344b CELLD r1=900e3 r0=10000e3
xl0b17c345 l0bl17 vdd x345 x345b CELLD r1=900e3 r0=10000e3
xl0b17c346 l0bl17 vdd x346 x346b CELLD r1=900e3 r0=10000e3
xl0b17c347 l0bl17 vdd x347 x347b CELLD r1=900e3 r0=10000e3
xl0b17c348 l0bl17 vdd x348 x348b CELLD r1=900e3 r0=10000e3
xl0b17c349 l0bl17 vdd x349 x349b CELLD r1=900e3 r0=10000e3
xl0b17c350 l0bl17 vdd x350 x350b CELLD r1=900e3 r0=10000e3
xl0b17c351 l0bl17 vdd x351 x351b CELLD r1=900e3 r0=10000e3
xl0b17c352 l0bl17 vdd x352 x352b CELLD r1=900e3 r0=10000e3
xl0b17c353 l0bl17 vdd x353 x353b CELLD r1=900e3 r0=10000e3
xl0b17c354 l0bl17 vdd x354 x354b CELLD r1=900e3 r0=10000e3
xl0b17c355 l0bl17 vdd x355 x355b CELLD r1=10000e3 r0=900e3
xl0b17c356 l0bl17 vdd x356 x356b CELLD r1=10000e3 r0=900e3
xl0b17c357 l0bl17 vdd x357 x357b CELLD r1=10000e3 r0=900e3
xl0b17c358 l0bl17 vdd x358 x358b CELLD r1=10000e3 r0=900e3
xl0b17c359 l0bl17 vdd x359 x359b CELLD r1=10000e3 r0=900e3
xl0b17c360 l0bl17 vdd x360 x360b CELLD r1=10000e3 r0=900e3
xl0b17c361 l0bl17 vdd x361 x361b CELLD r1=10000e3 r0=900e3
xl0b17c362 l0bl17 vdd x362 x362b CELLD r1=900e3 r0=10000e3
xl0b17c363 l0bl17 vdd x363 x363b CELLD r1=900e3 r0=10000e3
xl0b17c364 l0bl17 vdd x364 x364b CELLD r1=10000e3 r0=900e3
xl0b17c365 l0bl17 vdd x365 x365b CELLD r1=900e3 r0=10000e3
xl0b17c366 l0bl17 vdd x366 x366b CELLD r1=900e3 r0=10000e3
xl0b17c367 l0bl17 vdd x367 x367b CELLD r1=10000e3 r0=900e3
xl0b17c368 l0bl17 vdd x368 x368b CELLD r1=10000e3 r0=900e3
xl0b17c369 l0bl17 vdd x369 x369b CELLD r1=10000e3 r0=900e3
xl0b17c370 l0bl17 vdd x370 x370b CELLD r1=10000e3 r0=900e3
xl0b17c371 l0bl17 vdd x371 x371b CELLD r1=10000e3 r0=900e3
xl0b17c372 l0bl17 vdd x372 x372b CELLD r1=900e3 r0=10000e3
xl0b17c373 l0bl17 vdd x373 x373b CELLD r1=900e3 r0=10000e3
xl0b17c374 l0bl17 vdd x374 x374b CELLD r1=900e3 r0=10000e3
xl0b17c375 l0bl17 vdd x375 x375b CELLD r1=900e3 r0=10000e3
xl0b17c376 l0bl17 vdd x376 x376b CELLD r1=900e3 r0=10000e3
xl0b17c377 l0bl17 vdd x377 x377b CELLD r1=900e3 r0=10000e3
xl0b17c378 l0bl17 vdd x378 x378b CELLD r1=900e3 r0=10000e3
xl0b17c379 l0bl17 vdd x379 x379b CELLD r1=900e3 r0=10000e3
xl0b17c380 l0bl17 vdd x380 x380b CELLD r1=900e3 r0=10000e3
xl0b17c381 l0bl17 vdd x381 x381b CELLD r1=900e3 r0=10000e3
xl0b17c382 l0bl17 vdd x382 x382b CELLD r1=900e3 r0=10000e3
xl0b17c383 l0bl17 vdd x383 x383b CELLD r1=900e3 r0=10000e3
xl0b17c384 l0bl17 vdd x384 x384b CELLD r1=10000e3 r0=900e3
xl0b17c385 l0bl17 vdd x385 x385b CELLD r1=10000e3 r0=900e3
xl0b17c386 l0bl17 vdd x386 x386b CELLD r1=900e3 r0=10000e3
xl0b17c387 l0bl17 vdd x387 x387b CELLD r1=10000e3 r0=900e3
xl0b17c388 l0bl17 vdd x388 x388b CELLD r1=10000e3 r0=900e3
xl0b17c389 l0bl17 vdd x389 x389b CELLD r1=900e3 r0=10000e3
xl0b17c390 l0bl17 vdd x390 x390b CELLD r1=10000e3 r0=900e3
xl0b17c391 l0bl17 vdd x391 x391b CELLD r1=10000e3 r0=900e3
xl0b17c392 l0bl17 vdd x392 x392b CELLD r1=900e3 r0=10000e3
xl0b17c393 l0bl17 vdd x393 x393b CELLD r1=900e3 r0=10000e3
xl0b17c394 l0bl17 vdd x394 x394b CELLD r1=900e3 r0=10000e3
xl0b17c395 l0bl17 vdd x395 x395b CELLD r1=10000e3 r0=900e3
xl0b17c396 l0bl17 vdd x396 x396b CELLD r1=10000e3 r0=900e3
xl0b17c397 l0bl17 vdd x397 x397b CELLD r1=10000e3 r0=900e3
xl0b17c398 l0bl17 vdd x398 x398b CELLD r1=10000e3 r0=900e3
xl0b17c399 l0bl17 vdd x399 x399b CELLD r1=900e3 r0=10000e3
xl0b17c400 l0bl17 vdd x400 x400b CELLD r1=900e3 r0=10000e3
xl0b17c401 l0bl17 vdd x401 x401b CELLD r1=900e3 r0=10000e3
xl0b17c402 l0bl17 vdd x402 x402b CELLD r1=900e3 r0=10000e3
xl0b17c403 l0bl17 vdd x403 x403b CELLD r1=900e3 r0=10000e3
xl0b17c404 l0bl17 vdd x404 x404b CELLD r1=900e3 r0=10000e3
xl0b17c405 l0bl17 vdd x405 x405b CELLD r1=900e3 r0=10000e3
xl0b17c406 l0bl17 vdd x406 x406b CELLD r1=900e3 r0=10000e3
xl0b17c407 l0bl17 vdd x407 x407b CELLD r1=10000e3 r0=900e3
xl0b17c408 l0bl17 vdd x408 x408b CELLD r1=900e3 r0=10000e3
xl0b17c409 l0bl17 vdd x409 x409b CELLD r1=900e3 r0=10000e3
xl0b17c410 l0bl17 vdd x410 x410b CELLD r1=900e3 r0=10000e3
xl0b17c411 l0bl17 vdd x411 x411b CELLD r1=900e3 r0=10000e3
xl0b17c412 l0bl17 vdd x412 x412b CELLD r1=10000e3 r0=900e3
xl0b17c413 l0bl17 vdd x413 x413b CELLD r1=900e3 r0=10000e3
xl0b17c414 l0bl17 vdd x414 x414b CELLD r1=10000e3 r0=900e3
xl0b17c415 l0bl17 vdd x415 x415b CELLD r1=900e3 r0=10000e3
xl0b17c416 l0bl17 vdd x416 x416b CELLD r1=10000e3 r0=900e3
xl0b17c417 l0bl17 vdd x417 x417b CELLD r1=10000e3 r0=900e3
xl0b17c418 l0bl17 vdd x418 x418b CELLD r1=10000e3 r0=900e3
xl0b17c419 l0bl17 vdd x419 x419b CELLD r1=10000e3 r0=900e3
xl0b17c420 l0bl17 vdd x420 x420b CELLD r1=10000e3 r0=900e3
xl0b17c421 l0bl17 vdd x421 x421b CELLD r1=10000e3 r0=900e3
xl0b17c422 l0bl17 vdd x422 x422b CELLD r1=900e3 r0=10000e3
xl0b17c423 l0bl17 vdd x423 x423b CELLD r1=10000e3 r0=900e3
xl0b17c424 l0bl17 vdd x424 x424b CELLD r1=10000e3 r0=900e3
xl0b17c425 l0bl17 vdd x425 x425b CELLD r1=10000e3 r0=900e3
xl0b17c426 l0bl17 vdd x426 x426b CELLD r1=10000e3 r0=900e3
xl0b17c427 l0bl17 vdd x427 x427b CELLD r1=900e3 r0=10000e3
xl0b17c428 l0bl17 vdd x428 x428b CELLD r1=900e3 r0=10000e3
xl0b17c429 l0bl17 vdd x429 x429b CELLD r1=900e3 r0=10000e3
xl0b17c430 l0bl17 vdd x430 x430b CELLD r1=900e3 r0=10000e3
xl0b17c431 l0bl17 vdd x431 x431b CELLD r1=900e3 r0=10000e3
xl0b17c432 l0bl17 vdd x432 x432b CELLD r1=900e3 r0=10000e3
xl0b17c433 l0bl17 vdd x433 x433b CELLD r1=10000e3 r0=900e3
xl0b17c434 l0bl17 vdd x434 x434b CELLD r1=10000e3 r0=900e3
xl0b17c435 l0bl17 vdd x435 x435b CELLD r1=900e3 r0=10000e3
xl0b17c436 l0bl17 vdd x436 x436b CELLD r1=900e3 r0=10000e3
xl0b17c437 l0bl17 vdd x437 x437b CELLD r1=900e3 r0=10000e3
xl0b17c438 l0bl17 vdd x438 x438b CELLD r1=900e3 r0=10000e3
xl0b17c439 l0bl17 vdd x439 x439b CELLD r1=900e3 r0=10000e3
xl0b17c440 l0bl17 vdd x440 x440b CELLD r1=900e3 r0=10000e3
xl0b17c441 l0bl17 vdd x441 x441b CELLD r1=900e3 r0=10000e3
xl0b17c442 l0bl17 vdd x442 x442b CELLD r1=10000e3 r0=900e3
xl0b17c443 l0bl17 vdd x443 x443b CELLD r1=10000e3 r0=900e3
xl0b17c444 l0bl17 vdd x444 x444b CELLD r1=10000e3 r0=900e3
xl0b17c445 l0bl17 vdd x445 x445b CELLD r1=10000e3 r0=900e3
xl0b17c446 l0bl17 vdd x446 x446b CELLD r1=10000e3 r0=900e3
xl0b17c447 l0bl17 vdd x447 x447b CELLD r1=900e3 r0=10000e3
xl0b17c448 l0bl17 vdd x448 x448b CELLD r1=900e3 r0=10000e3
xl0b17c449 l0bl17 vdd x449 x449b CELLD r1=900e3 r0=10000e3
xl0b17c450 l0bl17 vdd x450 x450b CELLD r1=900e3 r0=10000e3
xl0b17c451 l0bl17 vdd x451 x451b CELLD r1=10000e3 r0=900e3
xl0b17c452 l0bl17 vdd x452 x452b CELLD r1=10000e3 r0=900e3
xl0b17c453 l0bl17 vdd x453 x453b CELLD r1=10000e3 r0=900e3
xl0b17c454 l0bl17 vdd x454 x454b CELLD r1=10000e3 r0=900e3
xl0b17c455 l0bl17 vdd x455 x455b CELLD r1=10000e3 r0=900e3
xl0b17c456 l0bl17 vdd x456 x456b CELLD r1=10000e3 r0=900e3
xl0b17c457 l0bl17 vdd x457 x457b CELLD r1=900e3 r0=10000e3
xl0b17c458 l0bl17 vdd x458 x458b CELLD r1=900e3 r0=10000e3
xl0b17c459 l0bl17 vdd x459 x459b CELLD r1=900e3 r0=10000e3
xl0b17c460 l0bl17 vdd x460 x460b CELLD r1=900e3 r0=10000e3
xl0b17c461 l0bl17 vdd x461 x461b CELLD r1=900e3 r0=10000e3
xl0b17c462 l0bl17 vdd x462 x462b CELLD r1=900e3 r0=10000e3
xl0b17c463 l0bl17 vdd x463 x463b CELLD r1=900e3 r0=10000e3
xl0b17c464 l0bl17 vdd x464 x464b CELLD r1=900e3 r0=10000e3
xl0b17c465 l0bl17 vdd x465 x465b CELLD r1=900e3 r0=10000e3
xl0b17c466 l0bl17 vdd x466 x466b CELLD r1=900e3 r0=10000e3
xl0b17c467 l0bl17 vdd x467 x467b CELLD r1=900e3 r0=10000e3
xl0b17c468 l0bl17 vdd x468 x468b CELLD r1=900e3 r0=10000e3
xl0b17c469 l0bl17 vdd x469 x469b CELLD r1=10000e3 r0=900e3
xl0b17c470 l0bl17 vdd x470 x470b CELLD r1=10000e3 r0=900e3
xl0b17c471 l0bl17 vdd x471 x471b CELLD r1=10000e3 r0=900e3
xl0b17c472 l0bl17 vdd x472 x472b CELLD r1=10000e3 r0=900e3
xl0b17c473 l0bl17 vdd x473 x473b CELLD r1=10000e3 r0=900e3
xl0b17c474 l0bl17 vdd x474 x474b CELLD r1=900e3 r0=10000e3
xl0b17c475 l0bl17 vdd x475 x475b CELLD r1=900e3 r0=10000e3
xl0b17c476 l0bl17 vdd x476 x476b CELLD r1=900e3 r0=10000e3
xl0b17c477 l0bl17 vdd x477 x477b CELLD r1=900e3 r0=10000e3
xl0b17c478 l0bl17 vdd x478 x478b CELLD r1=10000e3 r0=900e3
xl0b17c479 l0bl17 vdd x479 x479b CELLD r1=10000e3 r0=900e3
xl0b17c480 l0bl17 vdd x480 x480b CELLD r1=10000e3 r0=900e3
xl0b17c481 l0bl17 vdd x481 x481b CELLD r1=10000e3 r0=900e3
xl0b17c482 l0bl17 vdd x482 x482b CELLD r1=10000e3 r0=900e3
xl0b17c483 l0bl17 vdd x483 x483b CELLD r1=10000e3 r0=900e3
xl0b17c484 l0bl17 vdd x484 x484b CELLD r1=10000e3 r0=900e3
xl0b17c485 l0bl17 vdd x485 x485b CELLD r1=10000e3 r0=900e3
xl0b17c486 l0bl17 vdd x486 x486b CELLD r1=900e3 r0=10000e3
xl0b17c487 l0bl17 vdd x487 x487b CELLD r1=900e3 r0=10000e3
xl0b17c488 l0bl17 vdd x488 x488b CELLD r1=900e3 r0=10000e3
xl0b17c489 l0bl17 vdd x489 x489b CELLD r1=900e3 r0=10000e3
xl0b17c490 l0bl17 vdd x490 x490b CELLD r1=900e3 r0=10000e3
xl0b17c491 l0bl17 vdd x491 x491b CELLD r1=900e3 r0=10000e3
xl0b17c492 l0bl17 vdd x492 x492b CELLD r1=900e3 r0=10000e3
xl0b17c493 l0bl17 vdd x493 x493b CELLD r1=900e3 r0=10000e3
xl0b17c494 l0bl17 vdd x494 x494b CELLD r1=900e3 r0=10000e3
xl0b17c495 l0bl17 vdd x495 x495b CELLD r1=10000e3 r0=900e3
xl0b17c496 l0bl17 vdd x496 x496b CELLD r1=10000e3 r0=900e3
xl0b17c497 l0bl17 vdd x497 x497b CELLD r1=10000e3 r0=900e3
xl0b17c498 l0bl17 vdd x498 x498b CELLD r1=10000e3 r0=900e3
xl0b17c499 l0bl17 vdd x499 x499b CELLD r1=10000e3 r0=900e3
xl0b17c500 l0bl17 vdd x500 x500b CELLD r1=10000e3 r0=900e3
xl0b17c501 l0bl17 vdd x501 x501b CELLD r1=10000e3 r0=900e3
xl0b17c502 l0bl17 vdd x502 x502b CELLD r1=10000e3 r0=900e3
xl0b17c503 l0bl17 vdd x503 x503b CELLD r1=900e3 r0=10000e3
xl0b17c504 l0bl17 vdd x504 x504b CELLD r1=900e3 r0=10000e3
xl0b17c505 l0bl17 vdd x505 x505b CELLD r1=900e3 r0=10000e3
xl0b17c506 l0bl17 vdd x506 x506b CELLD r1=10000e3 r0=900e3
xl0b17c507 l0bl17 vdd x507 x507b CELLD r1=10000e3 r0=900e3
xl0b17c508 l0bl17 vdd x508 x508b CELLD r1=10000e3 r0=900e3
xl0b17c509 l0bl17 vdd x509 x509b CELLD r1=10000e3 r0=900e3
xl0b17c510 l0bl17 vdd x510 x510b CELLD r1=10000e3 r0=900e3
xl0b17c511 l0bl17 vdd x511 x511b CELLD r1=10000e3 r0=900e3
xl0b17c512 l0bl17 vdd x512 x512b CELLD r1=10000e3 r0=900e3
xl0b17c513 l0bl17 vdd x513 x513b CELLD r1=10000e3 r0=900e3
xl0b17c514 l0bl17 vdd x514 x514b CELLD r1=900e3 r0=10000e3
xl0b17c515 l0bl17 vdd x515 x515b CELLD r1=900e3 r0=10000e3
xl0b17c516 l0bl17 vdd x516 x516b CELLD r1=900e3 r0=10000e3
xl0b17c517 l0bl17 vdd x517 x517b CELLD r1=900e3 r0=10000e3
xl0b17c518 l0bl17 vdd x518 x518b CELLD r1=900e3 r0=10000e3
xl0b17c519 l0bl17 vdd x519 x519b CELLD r1=10000e3 r0=900e3
xl0b17c520 l0bl17 vdd x520 x520b CELLD r1=900e3 r0=10000e3
xl0b17c521 l0bl17 vdd x521 x521b CELLD r1=900e3 r0=10000e3
xl0b17c522 l0bl17 vdd x522 x522b CELLD r1=900e3 r0=10000e3
xl0b17c523 l0bl17 vdd x523 x523b CELLD r1=10000e3 r0=900e3
xl0b17c524 l0bl17 vdd x524 x524b CELLD r1=10000e3 r0=900e3
xl0b17c525 l0bl17 vdd x525 x525b CELLD r1=10000e3 r0=900e3
xl0b17c526 l0bl17 vdd x526 x526b CELLD r1=10000e3 r0=900e3
xl0b17c527 l0bl17 vdd x527 x527b CELLD r1=10000e3 r0=900e3
xl0b17c528 l0bl17 vdd x528 x528b CELLD r1=10000e3 r0=900e3
xl0b17c529 l0bl17 vdd x529 x529b CELLD r1=10000e3 r0=900e3
xl0b17c530 l0bl17 vdd x530 x530b CELLD r1=900e3 r0=10000e3
xl0b17c531 l0bl17 vdd x531 x531b CELLD r1=900e3 r0=10000e3
xl0b17c532 l0bl17 vdd x532 x532b CELLD r1=900e3 r0=10000e3
xl0b17c533 l0bl17 vdd x533 x533b CELLD r1=900e3 r0=10000e3
xl0b17c534 l0bl17 vdd x534 x534b CELLD r1=900e3 r0=10000e3
xl0b17c535 l0bl17 vdd x535 x535b CELLD r1=900e3 r0=10000e3
xl0b17c536 l0bl17 vdd x536 x536b CELLD r1=10000e3 r0=900e3
xl0b17c537 l0bl17 vdd x537 x537b CELLD r1=10000e3 r0=900e3
xl0b17c538 l0bl17 vdd x538 x538b CELLD r1=10000e3 r0=900e3
xl0b17c539 l0bl17 vdd x539 x539b CELLD r1=10000e3 r0=900e3
xl0b17c540 l0bl17 vdd x540 x540b CELLD r1=10000e3 r0=900e3
xl0b17c541 l0bl17 vdd x541 x541b CELLD r1=10000e3 r0=900e3
xl0b17c542 l0bl17 vdd x542 x542b CELLD r1=10000e3 r0=900e3
xl0b17c543 l0bl17 vdd x543 x543b CELLD r1=10000e3 r0=900e3
xl0b17c544 l0bl17 vdd x544 x544b CELLD r1=900e3 r0=10000e3
xl0b17c545 l0bl17 vdd x545 x545b CELLD r1=10000e3 r0=900e3
xl0b17c546 l0bl17 vdd x546 x546b CELLD r1=900e3 r0=10000e3
xl0b17c547 l0bl17 vdd x547 x547b CELLD r1=900e3 r0=10000e3
xl0b17c548 l0bl17 vdd x548 x548b CELLD r1=10000e3 r0=900e3
xl0b17c549 l0bl17 vdd x549 x549b CELLD r1=10000e3 r0=900e3
xl0b17c550 l0bl17 vdd x550 x550b CELLD r1=10000e3 r0=900e3
xl0b17c551 l0bl17 vdd x551 x551b CELLD r1=10000e3 r0=900e3
xl0b17c552 l0bl17 vdd x552 x552b CELLD r1=10000e3 r0=900e3
xl0b17c553 l0bl17 vdd x553 x553b CELLD r1=10000e3 r0=900e3
xl0b17c554 l0bl17 vdd x554 x554b CELLD r1=10000e3 r0=900e3
xl0b17c555 l0bl17 vdd x555 x555b CELLD r1=10000e3 r0=900e3
xl0b17c556 l0bl17 vdd x556 x556b CELLD r1=10000e3 r0=900e3
xl0b17c557 l0bl17 vdd x557 x557b CELLD r1=10000e3 r0=900e3
xl0b17c558 l0bl17 vdd x558 x558b CELLD r1=900e3 r0=10000e3
xl0b17c559 l0bl17 vdd x559 x559b CELLD r1=10000e3 r0=900e3
xl0b17c560 l0bl17 vdd x560 x560b CELLD r1=900e3 r0=10000e3
xl0b17c561 l0bl17 vdd x561 x561b CELLD r1=900e3 r0=10000e3
xl0b17c562 l0bl17 vdd x562 x562b CELLD r1=10000e3 r0=900e3
xl0b17c563 l0bl17 vdd x563 x563b CELLD r1=10000e3 r0=900e3
xl0b17c564 l0bl17 vdd x564 x564b CELLD r1=10000e3 r0=900e3
xl0b17c565 l0bl17 vdd x565 x565b CELLD r1=10000e3 r0=900e3
xl0b17c566 l0bl17 vdd x566 x566b CELLD r1=10000e3 r0=900e3
xl0b17c567 l0bl17 vdd x567 x567b CELLD r1=10000e3 r0=900e3
xl0b17c568 l0bl17 vdd x568 x568b CELLD r1=10000e3 r0=900e3
xl0b17c569 l0bl17 vdd x569 x569b CELLD r1=10000e3 r0=900e3
xl0b17c570 l0bl17 vdd x570 x570b CELLD r1=10000e3 r0=900e3
xl0b17c571 l0bl17 vdd x571 x571b CELLD r1=900e3 r0=10000e3
xl0b17c572 l0bl17 vdd x572 x572b CELLD r1=900e3 r0=10000e3
xl0b17c573 l0bl17 vdd x573 x573b CELLD r1=900e3 r0=10000e3
xl0b17c574 l0bl1